* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673769290314 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673769290310 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673769290313 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673769290311 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=6 EP=5 IP=10 FDC=3
X0 1 2 4 6 n18_CDNS_673769290310 $T=430 0 0 0 $X=110 $Y=-1130
X1 1 3 2 n18_CDNS_673769290313 $T=2660 100 0 0 $X=1960 $Y=-1130
X2 1 5 6 n18_CDNS_673769290311 $T=0 0 0 0 $X=-660 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_673769290312 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT DEC_AND CLK GND VDD A0 O0 A1 O1 A2 O2 A3 O3 A4 O4 A5 O5 A6 O6 A7 O7
** N=27 EP=19 IP=104 FDC=48
M0 VDD A0 5 VDD PM L=1.8e-07 W=8.8e-07 $X=-6315 $Y=4690 $D=4
M1 VDD A1 8 VDD PM L=1.8e-07 W=8.8e-07 $X=-1675 $Y=4690 $D=4
M2 VDD A2 11 VDD PM L=1.8e-07 W=8.8e-07 $X=2965 $Y=4690 $D=4
M3 VDD A3 14 VDD PM L=1.8e-07 W=8.8e-07 $X=7605 $Y=4690 $D=4
M4 VDD A4 17 VDD PM L=1.8e-07 W=8.8e-07 $X=12245 $Y=4690 $D=4
M5 VDD A5 20 VDD PM L=1.8e-07 W=8.8e-07 $X=16885 $Y=4690 $D=4
M6 VDD A6 23 VDD PM L=1.8e-07 W=8.8e-07 $X=21525 $Y=4690 $D=4
M7 VDD A7 26 VDD PM L=1.8e-07 W=8.8e-07 $X=26165 $Y=4690 $D=4
X8 VDD O0 5 p18_CDNS_673769290314 $T=-4375 5130 0 0 $X=-5285 $Y=4700
X9 VDD O1 8 p18_CDNS_673769290314 $T=265 5130 0 0 $X=-645 $Y=4700
X10 VDD O2 11 p18_CDNS_673769290314 $T=4905 5130 0 0 $X=3995 $Y=4700
X11 VDD O3 14 p18_CDNS_673769290314 $T=9545 5130 0 0 $X=8635 $Y=4700
X12 VDD O4 17 p18_CDNS_673769290314 $T=14185 5130 0 0 $X=13275 $Y=4700
X13 VDD O5 20 p18_CDNS_673769290314 $T=18825 5130 0 0 $X=17915 $Y=4700
X14 VDD O6 23 p18_CDNS_673769290314 $T=23465 5130 0 0 $X=22555 $Y=4700
X15 VDD O7 26 p18_CDNS_673769290314 $T=28105 5130 0 0 $X=27195 $Y=4700
X16 GND 5 O0 A0 CLK ICV_1 $T=-7035 -570 0 0 $X=-7695 $Y=-1700
X17 GND 8 O1 A1 CLK ICV_1 $T=-2395 -570 0 0 $X=-3055 $Y=-1700
X18 GND 11 O2 A2 CLK ICV_1 $T=2245 -570 0 0 $X=1585 $Y=-1700
X19 GND 14 O3 A3 CLK ICV_1 $T=6885 -570 0 0 $X=6225 $Y=-1700
X20 GND 17 O4 A4 CLK ICV_1 $T=11525 -570 0 0 $X=10865 $Y=-1700
X21 GND 20 O5 A5 CLK ICV_1 $T=16165 -570 0 0 $X=15505 $Y=-1700
X22 GND 23 O6 A6 CLK ICV_1 $T=20805 -570 0 0 $X=20145 $Y=-1700
X23 GND 26 O7 A7 CLK ICV_1 $T=25445 -570 0 0 $X=24785 $Y=-1700
X24 VDD 5 CLK p18_CDNS_673769290312 $T=-7035 4690 0 0 $X=-7945 $Y=4260
X25 VDD 8 CLK p18_CDNS_673769290312 $T=-2395 4690 0 0 $X=-3305 $Y=4260
X26 VDD 11 CLK p18_CDNS_673769290312 $T=2245 4690 0 0 $X=1335 $Y=4260
X27 VDD 14 CLK p18_CDNS_673769290312 $T=6885 4690 0 0 $X=5975 $Y=4260
X28 VDD 17 CLK p18_CDNS_673769290312 $T=11525 4690 0 0 $X=10615 $Y=4260
X29 VDD 20 CLK p18_CDNS_673769290312 $T=16165 4690 0 0 $X=15255 $Y=4260
X30 VDD 23 CLK p18_CDNS_673769290312 $T=20805 4690 0 0 $X=19895 $Y=4260
X31 VDD 26 CLK p18_CDNS_673769290312 $T=25445 4690 0 0 $X=24535 $Y=4260
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_673795915977 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159715 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 1 3 2 1 PM L=1.8e-07 W=3.3e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159716 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915976 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915979 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159710 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 5 6 n18_CDNS_673795915979 $T=0 -1660 0 0 $X=-660 $Y=-2010
X1 3 4 5 6 n18_CDNS_6737959159710 $T=0 0 0 0 $X=-660 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915972 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915973 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=16 FDC=4
X0 1 2 1 6 n18_CDNS_673795915972 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 1 3 7 n18_CDNS_673795915972 $T=2020 0 0 0 $X=1360 $Y=-1130
X2 1 2 4 8 n18_CDNS_673795915973 $T=0 2900 0 0 $X=-660 $Y=2550
X3 1 5 3 8 n18_CDNS_673795915973 $T=2020 2900 0 0 $X=1360 $Y=2550
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=8
X0 1 2 5 3 4 10 12 11 ICV_2 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 9 7 8 13 14 11 ICV_2 $T=4460 0 0 0 $X=3800 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159714 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4
** N=5 EP=4 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_6737959159714 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 1 4 p18_CDNS_6737959159714 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6
** N=7 EP=6 IP=10 FDC=4
X0 1 2 3 6 ICV_4 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 6 ICV_4 $T=4460 0 0 0 $X=3550 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_673795915974 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4
** N=5 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_673795915974 $T=-2020 0 0 0 $X=-2930 $Y=-1130
X1 1 3 2 p18_CDNS_673795915974 $T=0 0 0 0 $X=-910 $Y=-1130
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915978 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915975 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673795915978 $T=-2020 0 0 0 $X=-2720 $Y=-350
X1 1 3 2 n18_CDNS_673795915975 $T=0 0 0 0 $X=-700 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=8
X0 1 2 3 7 ICV_6 $T=-4460 0 0 0 $X=-7390 $Y=-1130
X1 1 4 5 8 ICV_6 $T=0 0 0 0 $X=-2930 $Y=-1130
X2 6 2 3 7 ICV_7 $T=-4460 1650 0 0 $X=-7180 $Y=1300
X3 6 4 5 8 ICV_7 $T=0 1650 0 0 $X=-2720 $Y=1300
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159712 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159711 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 n18_CDNS_6737959159712 $T=0 0 0 0 $X=-1520 $Y=-350
X1 3 1 2 n18_CDNS_6737959159711 $T=2020 0 0 0 $X=1360 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_9 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 4 5 ICV_9 $T=4460 0 0 0 $X=2940 $Y=-350
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159713 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3
** N=3 EP=3 IP=8 FDC=2
X0 1 1 2 3 p18_CDNS_6737959159713 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 3 1 2 p18_CDNS_6737959159713 $T=2020 0 0 0 $X=1070 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_11 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 4 5 ICV_11 $T=4460 0 0 0 $X=3510 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=20 FDC=16
X0 1 2 3 4 5 ICV_10 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 6 7 8 9 ICV_10 $T=8920 0 0 0 $X=7400 $Y=-350
X2 10 2 3 4 5 ICV_12 $T=0 1950 0 0 $X=-950 $Y=1420
X3 10 6 7 8 9 ICV_12 $T=8920 1950 0 0 $X=7970 $Y=1420
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=20 FDC=32
X0 1 3 4 5 6 7 8 9 10 2 ICV_13 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 11 12 13 14 15 16 17 18 2 ICV_13 $T=17840 0 0 0 $X=16320 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=34 EP=34 IP=36 FDC=64
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_14 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 2 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_14 $T=35680 0 0 0 $X=34160 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159723 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159726 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=3.52e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159725 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673795915970 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673795915970 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 3 2 n18_CDNS_673795915970 $T=1940 0 0 0 $X=1280 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159719 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_6737959159719 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 2 p18_CDNS_6737959159719 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159720 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159721 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4
** N=5 EP=4 IP=7 FDC=2
X0 1 3 5 p18_CDNS_6737959159720 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 2 4 5 p18_CDNS_6737959159721 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159717 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159722 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159724 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159718 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_6737959159717 $T=0 -1680 1 0 $X=-700 $Y=-2250
X1 1 3 5 n18_CDNS_6737959159717 $T=0 0 0 0 $X=-700 $Y=-1230
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_19 $T=0 0 0 0 $X=-700 $Y=-2250
X1 1 4 5 8 9 ICV_19 $T=2020 0 0 0 $X=1320 $Y=-2250
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_6737959159714 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 1 3 5 p18_CDNS_6737959159714 $T=0 2360 1 0 $X=-910 $Y=790
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_21 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 8 9 ICV_21 $T=2020 0 0 0 $X=1110 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 p18_CDNS_6737959159718 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 p18_CDNS_6737959159718 $T=0 3240 1 0 $X=-910 $Y=1230
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673795915970 $T=0 -1480 1 0 $X=-660 $Y=-2710
X1 1 3 5 n18_CDNS_673795915970 $T=0 0 0 0 $X=-660 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=4
X0 1 2 3 6 7 ICV_24 $T=0 0 0 0 $X=-660 $Y=-2710
X1 1 4 5 2 3 ICV_24 $T=1940 0 0 0 $X=1280 $Y=-2710
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7
** N=7 EP=7 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 7 ICV_17 $T=0 5000 1 0 $X=-910 $Y=2110
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_16 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 4 5 3 ICV_16 $T=3880 0 0 0 $X=3220 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=8
X0 1 2 3 4 5 10 ICV_27 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 7 8 9 5 ICV_27 $T=7760 0 0 0 $X=7100 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6
** N=7 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 3 ICV_17 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10
** N=11 EP=10 IP=14 FDC=8
X0 1 2 3 4 5 10 ICV_29 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 7 8 9 5 ICV_29 $T=7760 0 0 0 $X=6850 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=8
X0 1 2 4 3 5 10 11 ICV_26 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 8 7 9 4 5 ICV_26 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5
** N=6 EP=5 IP=10 FDC=3
X0 1 2 3 n18_CDNS_6737959159717 $T=0 0 0 0 $X=-700 $Y=-1230
X1 1 3 4 6 n18_CDNS_6737959159722 $T=-2230 -100 0 0 $X=-2550 $Y=-1230
X2 1 5 6 n18_CDNS_6737959159724 $T=-2660 -100 0 0 $X=-3320 $Y=-1230
.ENDS
***************************************
.SUBCKT p18_CDNS_673795915971 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159729 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 2 3 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6737959159728 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6737959159727 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT SRAM_8_16 A2 A1 A0 GND CLK MODE B0 INVB0 B1 INVB1 B2 INVB2 B3 INVB3 B4 INVB4 B5 INVB5 B6 INVB6
+ B7 INVB7 B8 INVB8 B9 INVB9 B10 INVB10 B11 INVB11 B12 INVB12 B13 INVB13 B14 INVB14 B15 INVB15 VDD CLKREG
+ ADD4 ADD3 SAEN ADD7 ADD6 ADD5 ADD2 ADD1 ADD0 O0 PCEN D0 O1 D1 O2 D2 O3 D3 O4 D4
+ O5 D5 O6 D6 O7 D7 O8 D8 O9 D9 O10 D10 O11 D11 O12 D12 O13 D13 O14 D14
+ O15 D15
** N=752 EP=82 IP=2653 FDC=1716
M0 GND A0 13 GND NM L=1.8e-07 W=2.2e-07 $X=-110655 $Y=-38680 $D=0
M1 GND 14 15 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-41920 $D=0
M2 15 13 GND GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-41120 $D=0
M3 18 12 GND GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-39100 $D=0
M4 GND 14 18 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-38300 $D=0
M5 GND A1 19 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-34680 $D=0
M6 GND A1 20 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-31060 $D=0
M7 GND 14 21 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-27440 $D=0
M8 GND 14 22 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-23820 $D=0
M9 GND A1 16 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-20200 $D=0
M10 GND A1 17 GND NM L=1.8e-07 W=2.2e-07 $X=-108935 $Y=-16580 $D=0
M11 194 25 GND GND NM L=1.8e-07 W=2.2e-07 $X=-95355 $Y=-1150 $D=0
M12 33 194 GND GND NM L=1.8e-07 W=2.2e-07 $X=-93335 $Y=-1150 $D=0
M13 198 196 GND GND NM L=1.8e-07 W=8.8e-07 $X=-92455 $Y=650 $D=0
M14 206 33 GND GND NM L=1.8e-07 W=8.8e-07 $X=-91355 $Y=-1710 $D=0
M15 216 206 GND GND NM L=1.8e-07 W=8.8e-07 $X=-89415 $Y=-1710 $D=0
M16 226 216 GND GND NM L=1.8e-07 W=8.8e-07 $X=-87475 $Y=-1710 $D=0
M17 236 226 GND GND NM L=1.8e-07 W=8.8e-07 $X=-85535 $Y=-1710 $D=0
M18 246 236 GND GND NM L=1.8e-07 W=8.8e-07 $X=-83595 $Y=-1710 $D=0
M19 257 246 GND GND NM L=1.8e-07 W=8.8e-07 $X=-81655 $Y=-1710 $D=0
M20 267 249 GND GND NM L=1.8e-07 W=8.8e-07 $X=-78875 $Y=650 $D=0
M21 276 33 708 GND NM L=1.8e-07 W=4.4e-07 $X=-77265 $Y=-1270 $D=0
M22 709 CLK GND GND NM L=1.8e-07 W=4.4e-07 $X=-74915 $Y=650 $D=0
M23 288 278 709 GND NM L=1.8e-07 W=4.4e-07 $X=-74485 $Y=650 $D=0
M24 290 280 710 GND NM L=1.8e-07 W=4.4e-07 $X=-72625 $Y=-60310 $D=0
M25 297 287 711 GND NM L=1.8e-07 W=4.4e-07 $X=-72625 $Y=-1270 $D=0
M26 298 290 GND GND NM L=1.8e-07 W=2.2e-07 $X=-70395 $Y=-60210 $D=0
M27 305 297 GND GND NM L=1.8e-07 W=2.2e-07 $X=-70395 $Y=-1150 $D=0
M28 40 298 GND GND NM L=1.8e-07 W=2.2e-07 $X=-68375 $Y=-60210 $D=0
M29 47 305 GND GND NM L=1.8e-07 W=2.2e-07 $X=-68375 $Y=-1150 $D=0
M30 50 1 GND GND NM L=1.8e-07 W=2.2e-07 $X=-66355 $Y=-60210 $D=0
M31 59 MODE 25 GND NM L=1.8e-07 W=4.4e-07 $X=-66235 $Y=650 $D=0
M32 24 36 58 GND NM L=1.8e-07 W=4.4e-07 $X=-65515 $Y=-62230 $D=0
M33 25 37 59 GND NM L=1.8e-07 W=4.4e-07 $X=-65515 $Y=650 $D=0
M34 58 38 GND GND NM L=1.8e-07 W=4.4e-07 $X=-63575 $Y=-62230 $D=0
M35 59 39 GND GND NM L=1.8e-07 W=4.4e-07 $X=-63575 $Y=650 $D=0
M36 GND 48 58 GND NM L=1.8e-07 W=4.4e-07 $X=-62855 $Y=-62230 $D=0
M37 GND 49 59 GND NM L=1.8e-07 W=4.4e-07 $X=-62855 $Y=650 $D=0
M38 ADD7 40 69 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-60310 $D=0
M39 ADD6 41 70 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-46990 $D=0
M40 ADD5 42 71 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-45070 $D=0
M41 ADD4 43 72 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-31750 $D=0
M42 ADD3 44 73 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-29830 $D=0
M43 ADD2 45 74 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-16510 $D=0
M44 ADD1 46 75 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-14590 $D=0
M45 ADD0 47 76 GND NM L=1.8e-07 W=4.4e-07 $X=-61635 $Y=-1270 $D=0
M46 76 57 GND GND NM L=1.8e-07 W=4.4e-07 $X=-59695 $Y=-1270 $D=0
M47 SAEN 311 GND GND NM L=1.8e-07 W=8.8e-07 $X=-58975 $Y=-62670 $D=0
M48 GND 61 69 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-60310 $D=0
M49 GND 62 70 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-46990 $D=0
M50 GND 63 71 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-45070 $D=0
M51 GND 64 72 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-31750 $D=0
M52 GND 65 73 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-29830 $D=0
M53 GND 66 74 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-16510 $D=0
M54 GND 67 75 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-14590 $D=0
M55 GND 68 76 GND NM L=1.8e-07 W=4.4e-07 $X=-58975 $Y=-1270 $D=0
M56 GND D0 78 GND NM L=1.8e-07 W=2.2e-07 $X=-54645 $Y=-67380 $D=0
M57 336 B0 326 GND NM L=1.8e-07 W=4.4e-07 $X=-54605 $Y=-58800 $D=0
M58 81 78 GND GND NM L=1.8e-07 W=2.2e-07 $X=-53845 $Y=-67380 $D=0
M59 GND D1 82 GND NM L=1.8e-07 W=2.2e-07 $X=-50185 $Y=-67380 $D=0
M60 360 B1 350 GND NM L=1.8e-07 W=4.4e-07 $X=-50145 $Y=-58800 $D=0
M61 85 82 GND GND NM L=1.8e-07 W=2.2e-07 $X=-49385 $Y=-67380 $D=0
M62 GND D2 86 GND NM L=1.8e-07 W=2.2e-07 $X=-45725 $Y=-67380 $D=0
M63 384 B2 374 GND NM L=1.8e-07 W=4.4e-07 $X=-45685 $Y=-58800 $D=0
M64 89 86 GND GND NM L=1.8e-07 W=2.2e-07 $X=-44925 $Y=-67380 $D=0
M65 GND D3 90 GND NM L=1.8e-07 W=2.2e-07 $X=-41265 $Y=-67380 $D=0
M66 408 B3 398 GND NM L=1.8e-07 W=4.4e-07 $X=-41225 $Y=-58800 $D=0
M67 93 90 GND GND NM L=1.8e-07 W=2.2e-07 $X=-40465 $Y=-67380 $D=0
M68 GND D4 94 GND NM L=1.8e-07 W=2.2e-07 $X=-36805 $Y=-67380 $D=0
M69 432 B4 422 GND NM L=1.8e-07 W=4.4e-07 $X=-36765 $Y=-58800 $D=0
M70 97 94 GND GND NM L=1.8e-07 W=2.2e-07 $X=-36005 $Y=-67380 $D=0
M71 GND D5 98 GND NM L=1.8e-07 W=2.2e-07 $X=-32345 $Y=-67380 $D=0
M72 456 B5 446 GND NM L=1.8e-07 W=4.4e-07 $X=-32305 $Y=-58800 $D=0
M73 101 98 GND GND NM L=1.8e-07 W=2.2e-07 $X=-31545 $Y=-67380 $D=0
M74 GND D6 102 GND NM L=1.8e-07 W=2.2e-07 $X=-27885 $Y=-67380 $D=0
M75 480 B6 470 GND NM L=1.8e-07 W=4.4e-07 $X=-27845 $Y=-58800 $D=0
M76 105 102 GND GND NM L=1.8e-07 W=2.2e-07 $X=-27085 $Y=-67380 $D=0
M77 GND D7 106 GND NM L=1.8e-07 W=2.2e-07 $X=-23425 $Y=-67380 $D=0
M78 504 B7 494 GND NM L=1.8e-07 W=4.4e-07 $X=-23385 $Y=-58800 $D=0
M79 109 106 GND GND NM L=1.8e-07 W=2.2e-07 $X=-22625 $Y=-67380 $D=0
M80 GND D8 110 GND NM L=1.8e-07 W=2.2e-07 $X=-18965 $Y=-67380 $D=0
M81 528 B8 518 GND NM L=1.8e-07 W=4.4e-07 $X=-18925 $Y=-58800 $D=0
M82 113 110 GND GND NM L=1.8e-07 W=2.2e-07 $X=-18165 $Y=-67380 $D=0
M83 GND D9 114 GND NM L=1.8e-07 W=2.2e-07 $X=-14505 $Y=-67380 $D=0
M84 552 B9 542 GND NM L=1.8e-07 W=4.4e-07 $X=-14465 $Y=-58800 $D=0
M85 117 114 GND GND NM L=1.8e-07 W=2.2e-07 $X=-13705 $Y=-67380 $D=0
M86 GND D10 118 GND NM L=1.8e-07 W=2.2e-07 $X=-10045 $Y=-67380 $D=0
M87 576 B10 566 GND NM L=1.8e-07 W=4.4e-07 $X=-10005 $Y=-58800 $D=0
M88 121 118 GND GND NM L=1.8e-07 W=2.2e-07 $X=-9245 $Y=-67380 $D=0
M89 GND D11 122 GND NM L=1.8e-07 W=2.2e-07 $X=-5585 $Y=-67380 $D=0
M90 600 B11 590 GND NM L=1.8e-07 W=4.4e-07 $X=-5545 $Y=-58800 $D=0
M91 125 122 GND GND NM L=1.8e-07 W=2.2e-07 $X=-4785 $Y=-67380 $D=0
M92 GND D12 126 GND NM L=1.8e-07 W=2.2e-07 $X=-1125 $Y=-67380 $D=0
M93 624 B12 614 GND NM L=1.8e-07 W=4.4e-07 $X=-1085 $Y=-58800 $D=0
M94 129 126 GND GND NM L=1.8e-07 W=2.2e-07 $X=-325 $Y=-67380 $D=0
M95 GND D13 130 GND NM L=1.8e-07 W=2.2e-07 $X=3335 $Y=-67380 $D=0
M96 648 B13 638 GND NM L=1.8e-07 W=4.4e-07 $X=3375 $Y=-58800 $D=0
M97 133 130 GND GND NM L=1.8e-07 W=2.2e-07 $X=4135 $Y=-67380 $D=0
M98 GND D14 134 GND NM L=1.8e-07 W=2.2e-07 $X=7795 $Y=-67380 $D=0
M99 672 B14 662 GND NM L=1.8e-07 W=4.4e-07 $X=7835 $Y=-58800 $D=0
M100 137 134 GND GND NM L=1.8e-07 W=2.2e-07 $X=8595 $Y=-67380 $D=0
M101 GND D15 138 GND NM L=1.8e-07 W=2.2e-07 $X=12255 $Y=-67380 $D=0
M102 696 B15 686 GND NM L=1.8e-07 W=4.4e-07 $X=12295 $Y=-58800 $D=0
M103 141 138 GND GND NM L=1.8e-07 W=2.2e-07 $X=13055 $Y=-67380 $D=0
M104 726 12 15 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-41980 $D=4
M105 VDD 13 727 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-41120 $D=4
M106 728 12 18 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-38360 $D=4
M107 729 14 728 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-37930 $D=4
M108 VDD A0 729 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-37500 $D=4
M109 730 12 19 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-34740 $D=4
M110 731 A1 730 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-34310 $D=4
M111 VDD 13 731 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-33880 $D=4
M112 VDD A0 732 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-30260 $D=4
M113 734 A1 733 VDD PM L=1.8e-07 W=1.32e-06 $X=-106765 $Y=-19830 $D=4
M114 176 15 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-48980 $D=4
M115 177 18 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-44340 $D=4
M116 178 19 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-39700 $D=4
M117 179 20 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-35060 $D=4
M118 180 21 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-30420 $D=4
M119 VDD 181 4 VDD PM L=1.8e-07 W=4.4e-07 $X=-103965 $Y=-27720 $D=4
M120 181 22 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-25780 $D=4
M121 VDD 182 3 VDD PM L=1.8e-07 W=4.4e-07 $X=-103965 $Y=-23080 $D=4
M122 182 16 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-21140 $D=4
M123 VDD CLK 182 VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-20420 $D=4
M124 183 17 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-16500 $D=4
M125 VDD CLK 183 VDD PM L=1.8e-07 W=8.8e-07 $X=-103965 $Y=-15780 $D=4
M126 VDD 26 269 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-55050 $D=4
M127 VDD 27 270 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-52690 $D=4
M128 VDD 28 271 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-39810 $D=4
M129 VDD 29 272 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-37450 $D=4
M130 VDD 30 273 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-24570 $D=4
M131 VDD 31 274 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-22210 $D=4
M132 VDD 32 275 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-9330 $D=4
M133 VDD 33 276 VDD PM L=1.8e-07 W=8.8e-07 $X=-76975 $Y=-6970 $D=4
M134 VDD 278 288 VDD PM L=1.8e-07 W=8.8e-07 $X=-74195 $Y=5910 $D=4
M135 VDD 280 290 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-55050 $D=4
M136 VDD 281 291 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-52690 $D=4
M137 VDD 282 292 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-39810 $D=4
M138 VDD 283 293 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-37450 $D=4
M139 VDD 284 294 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-24570 $D=4
M140 VDD 285 295 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-22210 $D=4
M141 VDD 286 296 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-9330 $D=4
M142 VDD 287 297 VDD PM L=1.8e-07 W=8.8e-07 $X=-72335 $Y=-6970 $D=4
M143 289 279 VDD VDD PM L=1.8e-07 W=1.76e-06 $X=-71455 $Y=-71170 $D=4
M144 38 GND VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-70235 $Y=-67930 $D=4
M145 307 306 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-67535 $Y=-69850 $D=4
M146 24 36 735 VDD PM L=1.8e-07 W=8.8e-07 $X=-65805 $Y=-67930 $D=4
M147 736 38 24 VDD PM L=1.8e-07 W=8.8e-07 $X=-65085 $Y=-67930 $D=4
M148 737 39 25 VDD PM L=1.8e-07 W=8.8e-07 $X=-65085 $Y=5910 $D=4
M149 VDD 307 308 VDD PM L=1.8e-07 W=8.8e-07 $X=-64835 $Y=-70290 $D=4
M150 VDD 48 736 VDD PM L=1.8e-07 W=8.8e-07 $X=-64655 $Y=-67930 $D=4
M151 VDD 49 737 VDD PM L=1.8e-07 W=8.8e-07 $X=-64655 $Y=5910 $D=4
M152 738 50 ADD7 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-55050 $D=4
M153 739 51 ADD6 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-52690 $D=4
M154 740 52 ADD5 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-39810 $D=4
M155 741 53 ADD4 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-37450 $D=4
M156 742 54 ADD3 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-24570 $D=4
M157 743 55 ADD2 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-22210 $D=4
M158 744 56 ADD1 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-9330 $D=4
M159 745 57 ADD0 VDD PM L=1.8e-07 W=8.8e-07 $X=-61205 $Y=-6970 $D=4
M160 VDD 61 738 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-55050 $D=4
M161 VDD 62 739 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-52690 $D=4
M162 VDD 63 740 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-39810 $D=4
M163 VDD 64 741 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-37450 $D=4
M164 VDD 65 742 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-24570 $D=4
M165 VDD 66 743 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-22210 $D=4
M166 VDD 67 744 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-9330 $D=4
M167 VDD 68 745 VDD PM L=1.8e-07 W=8.8e-07 $X=-60775 $Y=-6970 $D=4
M168 VDD D0 78 VDD PM L=1.8e-07 W=4.4e-07 $X=-54605 $Y=-65670 $D=4
M169 VDD 326 326 VDD PM L=1.8e-07 W=3.3e-06 $X=-54605 $Y=-56390 $D=4
M170 81 78 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-53885 $Y=-65670 $D=4
M171 VDD D1 82 VDD PM L=1.8e-07 W=4.4e-07 $X=-50145 $Y=-65670 $D=4
M172 VDD 350 350 VDD PM L=1.8e-07 W=3.3e-06 $X=-50145 $Y=-56390 $D=4
M173 85 82 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-49425 $Y=-65670 $D=4
M174 VDD D2 86 VDD PM L=1.8e-07 W=4.4e-07 $X=-45685 $Y=-65670 $D=4
M175 VDD 374 374 VDD PM L=1.8e-07 W=3.3e-06 $X=-45685 $Y=-56390 $D=4
M176 89 86 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-44965 $Y=-65670 $D=4
M177 VDD D3 90 VDD PM L=1.8e-07 W=4.4e-07 $X=-41225 $Y=-65670 $D=4
M178 VDD 398 398 VDD PM L=1.8e-07 W=3.3e-06 $X=-41225 $Y=-56390 $D=4
M179 93 90 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-40505 $Y=-65670 $D=4
M180 VDD D4 94 VDD PM L=1.8e-07 W=4.4e-07 $X=-36765 $Y=-65670 $D=4
M181 VDD 422 422 VDD PM L=1.8e-07 W=3.3e-06 $X=-36765 $Y=-56390 $D=4
M182 97 94 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-36045 $Y=-65670 $D=4
M183 VDD D5 98 VDD PM L=1.8e-07 W=4.4e-07 $X=-32305 $Y=-65670 $D=4
M184 VDD 446 446 VDD PM L=1.8e-07 W=3.3e-06 $X=-32305 $Y=-56390 $D=4
M185 101 98 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-31585 $Y=-65670 $D=4
M186 VDD D6 102 VDD PM L=1.8e-07 W=4.4e-07 $X=-27845 $Y=-65670 $D=4
M187 VDD 470 470 VDD PM L=1.8e-07 W=3.3e-06 $X=-27845 $Y=-56390 $D=4
M188 105 102 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-27125 $Y=-65670 $D=4
M189 VDD D7 106 VDD PM L=1.8e-07 W=4.4e-07 $X=-23385 $Y=-65670 $D=4
M190 VDD 494 494 VDD PM L=1.8e-07 W=3.3e-06 $X=-23385 $Y=-56390 $D=4
M191 109 106 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-22665 $Y=-65670 $D=4
M192 VDD D8 110 VDD PM L=1.8e-07 W=4.4e-07 $X=-18925 $Y=-65670 $D=4
M193 VDD 518 518 VDD PM L=1.8e-07 W=3.3e-06 $X=-18925 $Y=-56390 $D=4
M194 113 110 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-18205 $Y=-65670 $D=4
M195 VDD D9 114 VDD PM L=1.8e-07 W=4.4e-07 $X=-14465 $Y=-65670 $D=4
M196 VDD 542 542 VDD PM L=1.8e-07 W=3.3e-06 $X=-14465 $Y=-56390 $D=4
M197 117 114 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-13745 $Y=-65670 $D=4
M198 VDD D10 118 VDD PM L=1.8e-07 W=4.4e-07 $X=-10005 $Y=-65670 $D=4
M199 VDD 566 566 VDD PM L=1.8e-07 W=3.3e-06 $X=-10005 $Y=-56390 $D=4
M200 121 118 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-9285 $Y=-65670 $D=4
M201 VDD D11 122 VDD PM L=1.8e-07 W=4.4e-07 $X=-5545 $Y=-65670 $D=4
M202 VDD 590 590 VDD PM L=1.8e-07 W=3.3e-06 $X=-5545 $Y=-56390 $D=4
M203 125 122 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-4825 $Y=-65670 $D=4
M204 VDD D12 126 VDD PM L=1.8e-07 W=4.4e-07 $X=-1085 $Y=-65670 $D=4
M205 VDD 614 614 VDD PM L=1.8e-07 W=3.3e-06 $X=-1085 $Y=-56390 $D=4
M206 129 126 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-365 $Y=-65670 $D=4
M207 VDD D13 130 VDD PM L=1.8e-07 W=4.4e-07 $X=3375 $Y=-65670 $D=4
M208 VDD 638 638 VDD PM L=1.8e-07 W=3.3e-06 $X=3375 $Y=-56390 $D=4
M209 133 130 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=4095 $Y=-65670 $D=4
M210 VDD D14 134 VDD PM L=1.8e-07 W=4.4e-07 $X=7835 $Y=-65670 $D=4
M211 VDD 662 662 VDD PM L=1.8e-07 W=3.3e-06 $X=7835 $Y=-56390 $D=4
M212 137 134 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=8555 $Y=-65670 $D=4
M213 VDD D15 138 VDD PM L=1.8e-07 W=4.4e-07 $X=12295 $Y=-65670 $D=4
M214 VDD 686 686 VDD PM L=1.8e-07 W=3.3e-06 $X=12295 $Y=-56390 $D=4
M215 141 138 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=13015 $Y=-65670 $D=4
X216 GND 346 336 INVB0 n18_CDNS_673795915977 $T=-53705 -58800 1 180 $X=-54545 $Y=-59150
X217 GND 370 360 INVB1 n18_CDNS_673795915977 $T=-49245 -58800 1 180 $X=-50085 $Y=-59150
X218 GND 394 384 INVB2 n18_CDNS_673795915977 $T=-44785 -58800 1 180 $X=-45625 $Y=-59150
X219 GND 418 408 INVB3 n18_CDNS_673795915977 $T=-40325 -58800 1 180 $X=-41165 $Y=-59150
X220 GND 442 432 INVB4 n18_CDNS_673795915977 $T=-35865 -58800 1 180 $X=-36705 $Y=-59150
X221 GND 466 456 INVB5 n18_CDNS_673795915977 $T=-31405 -58800 1 180 $X=-32245 $Y=-59150
X222 GND 490 480 INVB6 n18_CDNS_673795915977 $T=-26945 -58800 1 180 $X=-27785 $Y=-59150
X223 GND 514 504 INVB7 n18_CDNS_673795915977 $T=-22485 -58800 1 180 $X=-23325 $Y=-59150
X224 GND 538 528 INVB8 n18_CDNS_673795915977 $T=-18025 -58800 1 180 $X=-18865 $Y=-59150
X225 GND 562 552 INVB9 n18_CDNS_673795915977 $T=-13565 -58800 1 180 $X=-14405 $Y=-59150
X226 GND 586 576 INVB10 n18_CDNS_673795915977 $T=-9105 -58800 1 180 $X=-9945 $Y=-59150
X227 GND 610 600 INVB11 n18_CDNS_673795915977 $T=-4645 -58800 1 180 $X=-5485 $Y=-59150
X228 GND 634 624 INVB12 n18_CDNS_673795915977 $T=-185 -58800 1 180 $X=-1025 $Y=-59150
X229 GND 658 648 INVB13 n18_CDNS_673795915977 $T=4275 -58800 1 180 $X=3435 $Y=-59150
X230 GND 682 672 INVB14 n18_CDNS_673795915977 $T=8735 -58800 1 180 $X=7895 $Y=-59150
X231 GND 706 696 INVB15 n18_CDNS_673795915977 $T=13195 -58800 1 180 $X=12355 $Y=-59150
X232 VDD 346 326 p18_CDNS_6737959159715 $T=-53705 -56390 1 180 $X=-54795 $Y=-56820
X233 VDD 370 350 p18_CDNS_6737959159715 $T=-49245 -56390 1 180 $X=-50335 $Y=-56820
X234 VDD 394 374 p18_CDNS_6737959159715 $T=-44785 -56390 1 180 $X=-45875 $Y=-56820
X235 VDD 418 398 p18_CDNS_6737959159715 $T=-40325 -56390 1 180 $X=-41415 $Y=-56820
X236 VDD 442 422 p18_CDNS_6737959159715 $T=-35865 -56390 1 180 $X=-36955 $Y=-56820
X237 VDD 466 446 p18_CDNS_6737959159715 $T=-31405 -56390 1 180 $X=-32495 $Y=-56820
X238 VDD 490 470 p18_CDNS_6737959159715 $T=-26945 -56390 1 180 $X=-28035 $Y=-56820
X239 VDD 514 494 p18_CDNS_6737959159715 $T=-22485 -56390 1 180 $X=-23575 $Y=-56820
X240 VDD 538 518 p18_CDNS_6737959159715 $T=-18025 -56390 1 180 $X=-19115 $Y=-56820
X241 VDD 562 542 p18_CDNS_6737959159715 $T=-13565 -56390 1 180 $X=-14655 $Y=-56820
X242 VDD 586 566 p18_CDNS_6737959159715 $T=-9105 -56390 1 180 $X=-10195 $Y=-56820
X243 VDD 610 590 p18_CDNS_6737959159715 $T=-4645 -56390 1 180 $X=-5735 $Y=-56820
X244 VDD 634 614 p18_CDNS_6737959159715 $T=-185 -56390 1 180 $X=-1275 $Y=-56820
X245 VDD 658 638 p18_CDNS_6737959159715 $T=4275 -56390 1 180 $X=3185 $Y=-56820
X246 VDD 682 662 p18_CDNS_6737959159715 $T=8735 -56390 1 180 $X=7645 $Y=-56820
X247 VDD 706 686 p18_CDNS_6737959159715 $T=13195 -56390 1 180 $X=12105 $Y=-56820
X248 B0 INVB0 PCEN VDD p18_CDNS_6737959159716 $T=-54375 -2720 0 270 $X=-54805 $Y=-3810
X249 B1 INVB1 PCEN VDD p18_CDNS_6737959159716 $T=-49915 -2720 0 270 $X=-50345 $Y=-3810
X250 B2 INVB2 PCEN VDD p18_CDNS_6737959159716 $T=-45455 -2720 0 270 $X=-45885 $Y=-3810
X251 B3 INVB3 PCEN VDD p18_CDNS_6737959159716 $T=-40995 -2720 0 270 $X=-41425 $Y=-3810
X252 B4 INVB4 PCEN VDD p18_CDNS_6737959159716 $T=-36535 -2720 0 270 $X=-36965 $Y=-3810
X253 B5 INVB5 PCEN VDD p18_CDNS_6737959159716 $T=-32075 -2720 0 270 $X=-32505 $Y=-3810
X254 B6 INVB6 PCEN VDD p18_CDNS_6737959159716 $T=-27615 -2720 0 270 $X=-28045 $Y=-3810
X255 B7 INVB7 PCEN VDD p18_CDNS_6737959159716 $T=-23155 -2720 0 270 $X=-23585 $Y=-3810
X256 B8 INVB8 PCEN VDD p18_CDNS_6737959159716 $T=-18695 -2720 0 270 $X=-19125 $Y=-3810
X257 B9 INVB9 PCEN VDD p18_CDNS_6737959159716 $T=-14235 -2720 0 270 $X=-14665 $Y=-3810
X258 B10 INVB10 PCEN VDD p18_CDNS_6737959159716 $T=-9775 -2720 0 270 $X=-10205 $Y=-3810
X259 B11 INVB11 PCEN VDD p18_CDNS_6737959159716 $T=-5315 -2720 0 270 $X=-5745 $Y=-3810
X260 B12 INVB12 PCEN VDD p18_CDNS_6737959159716 $T=-855 -2720 0 270 $X=-1285 $Y=-3810
X261 B13 INVB13 PCEN VDD p18_CDNS_6737959159716 $T=3605 -2720 0 270 $X=3175 $Y=-3810
X262 B14 INVB14 PCEN VDD p18_CDNS_6737959159716 $T=8065 -2720 0 270 $X=7635 $Y=-3810
X263 B15 INVB15 PCEN VDD p18_CDNS_6737959159716 $T=12525 -2720 0 270 $X=12095 $Y=-3810
X264 GND 336 SAEN n18_CDNS_673795915976 $T=-54595 -60430 1 90 $X=-54945 $Y=-61090
X265 GND 360 SAEN n18_CDNS_673795915976 $T=-50135 -60430 1 90 $X=-50485 $Y=-61090
X266 GND 384 SAEN n18_CDNS_673795915976 $T=-45675 -60430 1 90 $X=-46025 $Y=-61090
X267 GND 408 SAEN n18_CDNS_673795915976 $T=-41215 -60430 1 90 $X=-41565 $Y=-61090
X268 GND 432 SAEN n18_CDNS_673795915976 $T=-36755 -60430 1 90 $X=-37105 $Y=-61090
X269 GND 456 SAEN n18_CDNS_673795915976 $T=-32295 -60430 1 90 $X=-32645 $Y=-61090
X270 GND 480 SAEN n18_CDNS_673795915976 $T=-27835 -60430 1 90 $X=-28185 $Y=-61090
X271 GND 504 SAEN n18_CDNS_673795915976 $T=-23375 -60430 1 90 $X=-23725 $Y=-61090
X272 GND 528 SAEN n18_CDNS_673795915976 $T=-18915 -60430 1 90 $X=-19265 $Y=-61090
X273 GND 552 SAEN n18_CDNS_673795915976 $T=-14455 -60430 1 90 $X=-14805 $Y=-61090
X274 GND 576 SAEN n18_CDNS_673795915976 $T=-9995 -60430 1 90 $X=-10345 $Y=-61090
X275 GND 600 SAEN n18_CDNS_673795915976 $T=-5535 -60430 1 90 $X=-5885 $Y=-61090
X276 GND 624 SAEN n18_CDNS_673795915976 $T=-1075 -60430 1 90 $X=-1425 $Y=-61090
X277 GND 648 SAEN n18_CDNS_673795915976 $T=3385 -60430 1 90 $X=3035 $Y=-61090
X278 GND 672 SAEN n18_CDNS_673795915976 $T=7845 -60430 1 90 $X=7495 $Y=-61090
X279 GND 696 SAEN n18_CDNS_673795915976 $T=12305 -60430 1 90 $X=11955 $Y=-61090
X280 INVB0 338 B0 327 ADD7 GND ICV_1 $T=-54765 -50860 0 90 $X=-55555 $Y=-51520
X281 INVB0 339 B0 328 ADD6 GND ICV_1 $T=-54765 -44820 0 90 $X=-55555 $Y=-45480
X282 INVB0 340 B0 329 ADD5 GND ICV_1 $T=-54765 -38780 0 90 $X=-55555 $Y=-39440
X283 INVB0 341 B0 330 ADD4 GND ICV_1 $T=-54765 -32740 0 90 $X=-55555 $Y=-33400
X284 INVB0 342 B0 331 ADD3 GND ICV_1 $T=-54765 -26700 0 90 $X=-55555 $Y=-27360
X285 INVB0 343 B0 332 ADD2 GND ICV_1 $T=-54765 -20660 0 90 $X=-55555 $Y=-21320
X286 INVB0 344 B0 333 ADD1 GND ICV_1 $T=-54765 -14620 0 90 $X=-55555 $Y=-15280
X287 INVB0 345 B0 334 ADD0 GND ICV_1 $T=-54765 -8580 0 90 $X=-55555 $Y=-9240
X288 INVB1 362 B1 351 ADD7 GND ICV_1 $T=-50305 -50860 0 90 $X=-51095 $Y=-51520
X289 INVB1 363 B1 352 ADD6 GND ICV_1 $T=-50305 -44820 0 90 $X=-51095 $Y=-45480
X290 INVB1 364 B1 353 ADD5 GND ICV_1 $T=-50305 -38780 0 90 $X=-51095 $Y=-39440
X291 INVB1 365 B1 354 ADD4 GND ICV_1 $T=-50305 -32740 0 90 $X=-51095 $Y=-33400
X292 INVB1 366 B1 355 ADD3 GND ICV_1 $T=-50305 -26700 0 90 $X=-51095 $Y=-27360
X293 INVB1 367 B1 356 ADD2 GND ICV_1 $T=-50305 -20660 0 90 $X=-51095 $Y=-21320
X294 INVB1 368 B1 357 ADD1 GND ICV_1 $T=-50305 -14620 0 90 $X=-51095 $Y=-15280
X295 INVB1 369 B1 358 ADD0 GND ICV_1 $T=-50305 -8580 0 90 $X=-51095 $Y=-9240
X296 INVB2 386 B2 375 ADD7 GND ICV_1 $T=-45845 -50860 0 90 $X=-46635 $Y=-51520
X297 INVB2 387 B2 376 ADD6 GND ICV_1 $T=-45845 -44820 0 90 $X=-46635 $Y=-45480
X298 INVB2 388 B2 377 ADD5 GND ICV_1 $T=-45845 -38780 0 90 $X=-46635 $Y=-39440
X299 INVB2 389 B2 378 ADD4 GND ICV_1 $T=-45845 -32740 0 90 $X=-46635 $Y=-33400
X300 INVB2 390 B2 379 ADD3 GND ICV_1 $T=-45845 -26700 0 90 $X=-46635 $Y=-27360
X301 INVB2 391 B2 380 ADD2 GND ICV_1 $T=-45845 -20660 0 90 $X=-46635 $Y=-21320
X302 INVB2 392 B2 381 ADD1 GND ICV_1 $T=-45845 -14620 0 90 $X=-46635 $Y=-15280
X303 INVB2 393 B2 382 ADD0 GND ICV_1 $T=-45845 -8580 0 90 $X=-46635 $Y=-9240
X304 INVB3 410 B3 399 ADD7 GND ICV_1 $T=-41385 -50860 0 90 $X=-42175 $Y=-51520
X305 INVB3 411 B3 400 ADD6 GND ICV_1 $T=-41385 -44820 0 90 $X=-42175 $Y=-45480
X306 INVB3 412 B3 401 ADD5 GND ICV_1 $T=-41385 -38780 0 90 $X=-42175 $Y=-39440
X307 INVB3 413 B3 402 ADD4 GND ICV_1 $T=-41385 -32740 0 90 $X=-42175 $Y=-33400
X308 INVB3 414 B3 403 ADD3 GND ICV_1 $T=-41385 -26700 0 90 $X=-42175 $Y=-27360
X309 INVB3 415 B3 404 ADD2 GND ICV_1 $T=-41385 -20660 0 90 $X=-42175 $Y=-21320
X310 INVB3 416 B3 405 ADD1 GND ICV_1 $T=-41385 -14620 0 90 $X=-42175 $Y=-15280
X311 INVB3 417 B3 406 ADD0 GND ICV_1 $T=-41385 -8580 0 90 $X=-42175 $Y=-9240
X312 INVB4 434 B4 423 ADD7 GND ICV_1 $T=-36925 -50860 0 90 $X=-37715 $Y=-51520
X313 INVB4 435 B4 424 ADD6 GND ICV_1 $T=-36925 -44820 0 90 $X=-37715 $Y=-45480
X314 INVB4 436 B4 425 ADD5 GND ICV_1 $T=-36925 -38780 0 90 $X=-37715 $Y=-39440
X315 INVB4 437 B4 426 ADD4 GND ICV_1 $T=-36925 -32740 0 90 $X=-37715 $Y=-33400
X316 INVB4 438 B4 427 ADD3 GND ICV_1 $T=-36925 -26700 0 90 $X=-37715 $Y=-27360
X317 INVB4 439 B4 428 ADD2 GND ICV_1 $T=-36925 -20660 0 90 $X=-37715 $Y=-21320
X318 INVB4 440 B4 429 ADD1 GND ICV_1 $T=-36925 -14620 0 90 $X=-37715 $Y=-15280
X319 INVB4 441 B4 430 ADD0 GND ICV_1 $T=-36925 -8580 0 90 $X=-37715 $Y=-9240
X320 INVB5 458 B5 447 ADD7 GND ICV_1 $T=-32465 -50860 0 90 $X=-33255 $Y=-51520
X321 INVB5 459 B5 448 ADD6 GND ICV_1 $T=-32465 -44820 0 90 $X=-33255 $Y=-45480
X322 INVB5 460 B5 449 ADD5 GND ICV_1 $T=-32465 -38780 0 90 $X=-33255 $Y=-39440
X323 INVB5 461 B5 450 ADD4 GND ICV_1 $T=-32465 -32740 0 90 $X=-33255 $Y=-33400
X324 INVB5 462 B5 451 ADD3 GND ICV_1 $T=-32465 -26700 0 90 $X=-33255 $Y=-27360
X325 INVB5 463 B5 452 ADD2 GND ICV_1 $T=-32465 -20660 0 90 $X=-33255 $Y=-21320
X326 INVB5 464 B5 453 ADD1 GND ICV_1 $T=-32465 -14620 0 90 $X=-33255 $Y=-15280
X327 INVB5 465 B5 454 ADD0 GND ICV_1 $T=-32465 -8580 0 90 $X=-33255 $Y=-9240
X328 INVB6 482 B6 471 ADD7 GND ICV_1 $T=-28005 -50860 0 90 $X=-28795 $Y=-51520
X329 INVB6 483 B6 472 ADD6 GND ICV_1 $T=-28005 -44820 0 90 $X=-28795 $Y=-45480
X330 INVB6 484 B6 473 ADD5 GND ICV_1 $T=-28005 -38780 0 90 $X=-28795 $Y=-39440
X331 INVB6 485 B6 474 ADD4 GND ICV_1 $T=-28005 -32740 0 90 $X=-28795 $Y=-33400
X332 INVB6 486 B6 475 ADD3 GND ICV_1 $T=-28005 -26700 0 90 $X=-28795 $Y=-27360
X333 INVB6 487 B6 476 ADD2 GND ICV_1 $T=-28005 -20660 0 90 $X=-28795 $Y=-21320
X334 INVB6 488 B6 477 ADD1 GND ICV_1 $T=-28005 -14620 0 90 $X=-28795 $Y=-15280
X335 INVB6 489 B6 478 ADD0 GND ICV_1 $T=-28005 -8580 0 90 $X=-28795 $Y=-9240
X336 INVB7 506 B7 495 ADD7 GND ICV_1 $T=-23545 -50860 0 90 $X=-24335 $Y=-51520
X337 INVB7 507 B7 496 ADD6 GND ICV_1 $T=-23545 -44820 0 90 $X=-24335 $Y=-45480
X338 INVB7 508 B7 497 ADD5 GND ICV_1 $T=-23545 -38780 0 90 $X=-24335 $Y=-39440
X339 INVB7 509 B7 498 ADD4 GND ICV_1 $T=-23545 -32740 0 90 $X=-24335 $Y=-33400
X340 INVB7 510 B7 499 ADD3 GND ICV_1 $T=-23545 -26700 0 90 $X=-24335 $Y=-27360
X341 INVB7 511 B7 500 ADD2 GND ICV_1 $T=-23545 -20660 0 90 $X=-24335 $Y=-21320
X342 INVB7 512 B7 501 ADD1 GND ICV_1 $T=-23545 -14620 0 90 $X=-24335 $Y=-15280
X343 INVB7 513 B7 502 ADD0 GND ICV_1 $T=-23545 -8580 0 90 $X=-24335 $Y=-9240
X344 INVB8 530 B8 519 ADD7 GND ICV_1 $T=-19085 -50860 0 90 $X=-19875 $Y=-51520
X345 INVB8 531 B8 520 ADD6 GND ICV_1 $T=-19085 -44820 0 90 $X=-19875 $Y=-45480
X346 INVB8 532 B8 521 ADD5 GND ICV_1 $T=-19085 -38780 0 90 $X=-19875 $Y=-39440
X347 INVB8 533 B8 522 ADD4 GND ICV_1 $T=-19085 -32740 0 90 $X=-19875 $Y=-33400
X348 INVB8 534 B8 523 ADD3 GND ICV_1 $T=-19085 -26700 0 90 $X=-19875 $Y=-27360
X349 INVB8 535 B8 524 ADD2 GND ICV_1 $T=-19085 -20660 0 90 $X=-19875 $Y=-21320
X350 INVB8 536 B8 525 ADD1 GND ICV_1 $T=-19085 -14620 0 90 $X=-19875 $Y=-15280
X351 INVB8 537 B8 526 ADD0 GND ICV_1 $T=-19085 -8580 0 90 $X=-19875 $Y=-9240
X352 INVB9 554 B9 543 ADD7 GND ICV_1 $T=-14625 -50860 0 90 $X=-15415 $Y=-51520
X353 INVB9 555 B9 544 ADD6 GND ICV_1 $T=-14625 -44820 0 90 $X=-15415 $Y=-45480
X354 INVB9 556 B9 545 ADD5 GND ICV_1 $T=-14625 -38780 0 90 $X=-15415 $Y=-39440
X355 INVB9 557 B9 546 ADD4 GND ICV_1 $T=-14625 -32740 0 90 $X=-15415 $Y=-33400
X356 INVB9 558 B9 547 ADD3 GND ICV_1 $T=-14625 -26700 0 90 $X=-15415 $Y=-27360
X357 INVB9 559 B9 548 ADD2 GND ICV_1 $T=-14625 -20660 0 90 $X=-15415 $Y=-21320
X358 INVB9 560 B9 549 ADD1 GND ICV_1 $T=-14625 -14620 0 90 $X=-15415 $Y=-15280
X359 INVB9 561 B9 550 ADD0 GND ICV_1 $T=-14625 -8580 0 90 $X=-15415 $Y=-9240
X360 INVB10 578 B10 567 ADD7 GND ICV_1 $T=-10165 -50860 0 90 $X=-10955 $Y=-51520
X361 INVB10 579 B10 568 ADD6 GND ICV_1 $T=-10165 -44820 0 90 $X=-10955 $Y=-45480
X362 INVB10 580 B10 569 ADD5 GND ICV_1 $T=-10165 -38780 0 90 $X=-10955 $Y=-39440
X363 INVB10 581 B10 570 ADD4 GND ICV_1 $T=-10165 -32740 0 90 $X=-10955 $Y=-33400
X364 INVB10 582 B10 571 ADD3 GND ICV_1 $T=-10165 -26700 0 90 $X=-10955 $Y=-27360
X365 INVB10 583 B10 572 ADD2 GND ICV_1 $T=-10165 -20660 0 90 $X=-10955 $Y=-21320
X366 INVB10 584 B10 573 ADD1 GND ICV_1 $T=-10165 -14620 0 90 $X=-10955 $Y=-15280
X367 INVB10 585 B10 574 ADD0 GND ICV_1 $T=-10165 -8580 0 90 $X=-10955 $Y=-9240
X368 INVB11 602 B11 591 ADD7 GND ICV_1 $T=-5705 -50860 0 90 $X=-6495 $Y=-51520
X369 INVB11 603 B11 592 ADD6 GND ICV_1 $T=-5705 -44820 0 90 $X=-6495 $Y=-45480
X370 INVB11 604 B11 593 ADD5 GND ICV_1 $T=-5705 -38780 0 90 $X=-6495 $Y=-39440
X371 INVB11 605 B11 594 ADD4 GND ICV_1 $T=-5705 -32740 0 90 $X=-6495 $Y=-33400
X372 INVB11 606 B11 595 ADD3 GND ICV_1 $T=-5705 -26700 0 90 $X=-6495 $Y=-27360
X373 INVB11 607 B11 596 ADD2 GND ICV_1 $T=-5705 -20660 0 90 $X=-6495 $Y=-21320
X374 INVB11 608 B11 597 ADD1 GND ICV_1 $T=-5705 -14620 0 90 $X=-6495 $Y=-15280
X375 INVB11 609 B11 598 ADD0 GND ICV_1 $T=-5705 -8580 0 90 $X=-6495 $Y=-9240
X376 INVB12 626 B12 615 ADD7 GND ICV_1 $T=-1245 -50860 0 90 $X=-2035 $Y=-51520
X377 INVB12 627 B12 616 ADD6 GND ICV_1 $T=-1245 -44820 0 90 $X=-2035 $Y=-45480
X378 INVB12 628 B12 617 ADD5 GND ICV_1 $T=-1245 -38780 0 90 $X=-2035 $Y=-39440
X379 INVB12 629 B12 618 ADD4 GND ICV_1 $T=-1245 -32740 0 90 $X=-2035 $Y=-33400
X380 INVB12 630 B12 619 ADD3 GND ICV_1 $T=-1245 -26700 0 90 $X=-2035 $Y=-27360
X381 INVB12 631 B12 620 ADD2 GND ICV_1 $T=-1245 -20660 0 90 $X=-2035 $Y=-21320
X382 INVB12 632 B12 621 ADD1 GND ICV_1 $T=-1245 -14620 0 90 $X=-2035 $Y=-15280
X383 INVB12 633 B12 622 ADD0 GND ICV_1 $T=-1245 -8580 0 90 $X=-2035 $Y=-9240
X384 INVB13 650 B13 639 ADD7 GND ICV_1 $T=3215 -50860 0 90 $X=2425 $Y=-51520
X385 INVB13 651 B13 640 ADD6 GND ICV_1 $T=3215 -44820 0 90 $X=2425 $Y=-45480
X386 INVB13 652 B13 641 ADD5 GND ICV_1 $T=3215 -38780 0 90 $X=2425 $Y=-39440
X387 INVB13 653 B13 642 ADD4 GND ICV_1 $T=3215 -32740 0 90 $X=2425 $Y=-33400
X388 INVB13 654 B13 643 ADD3 GND ICV_1 $T=3215 -26700 0 90 $X=2425 $Y=-27360
X389 INVB13 655 B13 644 ADD2 GND ICV_1 $T=3215 -20660 0 90 $X=2425 $Y=-21320
X390 INVB13 656 B13 645 ADD1 GND ICV_1 $T=3215 -14620 0 90 $X=2425 $Y=-15280
X391 INVB13 657 B13 646 ADD0 GND ICV_1 $T=3215 -8580 0 90 $X=2425 $Y=-9240
X392 INVB14 674 B14 663 ADD7 GND ICV_1 $T=7675 -50860 0 90 $X=6885 $Y=-51520
X393 INVB14 675 B14 664 ADD6 GND ICV_1 $T=7675 -44820 0 90 $X=6885 $Y=-45480
X394 INVB14 676 B14 665 ADD5 GND ICV_1 $T=7675 -38780 0 90 $X=6885 $Y=-39440
X395 INVB14 677 B14 666 ADD4 GND ICV_1 $T=7675 -32740 0 90 $X=6885 $Y=-33400
X396 INVB14 678 B14 667 ADD3 GND ICV_1 $T=7675 -26700 0 90 $X=6885 $Y=-27360
X397 INVB14 679 B14 668 ADD2 GND ICV_1 $T=7675 -20660 0 90 $X=6885 $Y=-21320
X398 INVB14 680 B14 669 ADD1 GND ICV_1 $T=7675 -14620 0 90 $X=6885 $Y=-15280
X399 INVB14 681 B14 670 ADD0 GND ICV_1 $T=7675 -8580 0 90 $X=6885 $Y=-9240
X400 INVB15 698 B15 687 ADD7 GND ICV_1 $T=12135 -50860 0 90 $X=11345 $Y=-51520
X401 INVB15 699 B15 688 ADD6 GND ICV_1 $T=12135 -44820 0 90 $X=11345 $Y=-45480
X402 INVB15 700 B15 689 ADD5 GND ICV_1 $T=12135 -38780 0 90 $X=11345 $Y=-39440
X403 INVB15 701 B15 690 ADD4 GND ICV_1 $T=12135 -32740 0 90 $X=11345 $Y=-33400
X404 INVB15 702 B15 691 ADD3 GND ICV_1 $T=12135 -26700 0 90 $X=11345 $Y=-27360
X405 INVB15 703 B15 692 ADD2 GND ICV_1 $T=12135 -20660 0 90 $X=11345 $Y=-21320
X406 INVB15 704 B15 693 ADD1 GND ICV_1 $T=12135 -14620 0 90 $X=11345 $Y=-15280
X407 INVB15 705 B15 694 ADD0 GND ICV_1 $T=12135 -8580 0 90 $X=11345 $Y=-9240
X408 GND 324 B0 INVB0 347 349 B1 INVB1 371 78 MODE 81 82 85 ICV_3 $T=-55255 -73530 0 0 $X=-55915 $Y=-74660
X409 GND 373 B2 INVB2 395 397 B3 INVB3 419 86 MODE 89 90 93 ICV_3 $T=-46335 -73530 0 0 $X=-46995 $Y=-74660
X410 GND 421 B4 INVB4 443 445 B5 INVB5 467 94 MODE 97 98 101 ICV_3 $T=-37415 -73530 0 0 $X=-38075 $Y=-74660
X411 GND 469 B6 INVB6 491 493 B7 INVB7 515 102 MODE 105 106 109 ICV_3 $T=-28495 -73530 0 0 $X=-29155 $Y=-74660
X412 GND 517 B8 INVB8 539 541 B9 INVB9 563 110 MODE 113 114 117 ICV_3 $T=-19575 -73530 0 0 $X=-20235 $Y=-74660
X413 GND 565 B10 INVB10 587 589 B11 INVB11 611 118 MODE 121 122 125 ICV_3 $T=-10655 -73530 0 0 $X=-11315 $Y=-74660
X414 GND 613 B12 INVB12 635 637 B13 INVB13 659 126 MODE 129 130 133 ICV_3 $T=-1735 -73530 0 0 $X=-2395 $Y=-74660
X415 GND 661 B14 INVB14 683 685 B15 INVB15 707 134 MODE 137 138 141 ICV_3 $T=7185 -73530 0 0 $X=6525 $Y=-74660
X416 VDD VDD 12 A2 p18_CDNS_6737959159714 $T=-113970 -42540 1 270 $X=-115540 $Y=-43630
X417 VDD VDD 14 A1 p18_CDNS_6737959159714 $T=-113970 -40520 1 270 $X=-115540 $Y=-41610
X418 VDD VDD 13 A0 p18_CDNS_6737959159714 $T=-113970 -38500 1 270 $X=-115540 $Y=-39590
X419 VDD VDD 1 176 p18_CDNS_6737959159714 $T=-103525 -50740 1 270 $X=-105095 $Y=-51830
X420 VDD VDD 6 177 p18_CDNS_6737959159714 $T=-103525 -46100 1 270 $X=-105095 $Y=-47190
X421 VDD VDD 5 178 p18_CDNS_6737959159714 $T=-103525 -41460 1 270 $X=-105095 $Y=-42550
X422 VDD VDD 7 179 p18_CDNS_6737959159714 $T=-103525 -36820 1 270 $X=-105095 $Y=-37910
X423 VDD VDD 8 180 p18_CDNS_6737959159714 $T=-103525 -32180 1 270 $X=-105095 $Y=-33270
X424 VDD VDD 2 183 p18_CDNS_6737959159714 $T=-103525 -18260 1 270 $X=-105095 $Y=-19350
X425 VDD VDD 278 267 p18_CDNS_6737959159714 $T=-76895 6350 0 0 $X=-77805 $Y=5920
X426 VDD VDD 36 34 p18_CDNS_6737959159714 $T=-72255 -67490 1 0 $X=-73165 $Y=-69060
X427 VDD VDD 37 288 p18_CDNS_6737959159714 $T=-72255 6350 0 0 $X=-73165 $Y=5920
X428 VDD VDD 39 VDD p18_CDNS_6737959159714 $T=-70235 6350 0 0 $X=-71145 $Y=5920
X429 VDD VDD 48 MODE p18_CDNS_6737959159714 $T=-68215 -67490 1 0 $X=-69125 $Y=-69060
X430 VDD VDD 49 MODE p18_CDNS_6737959159714 $T=-68215 6350 0 0 $X=-69125 $Y=5920
X431 VDD VDD 309 308 p18_CDNS_6737959159714 $T=-62895 -69850 0 0 $X=-63805 $Y=-70280
X432 VDD B0 INVB0 B1 INVB1 PCEN ICV_5 $T=-55215 -1270 0 0 $X=-56125 $Y=-1700
X433 VDD B2 INVB2 B3 INVB3 PCEN ICV_5 $T=-46295 -1270 0 0 $X=-47205 $Y=-1700
X434 VDD B4 INVB4 B5 INVB5 PCEN ICV_5 $T=-37375 -1270 0 0 $X=-38285 $Y=-1700
X435 VDD B6 INVB6 B7 INVB7 PCEN ICV_5 $T=-28455 -1270 0 0 $X=-29365 $Y=-1700
X436 VDD B8 INVB8 B9 INVB9 PCEN ICV_5 $T=-19535 -1270 0 0 $X=-20445 $Y=-1700
X437 VDD B10 INVB10 B11 INVB11 PCEN ICV_5 $T=-10615 -1270 0 0 $X=-11525 $Y=-1700
X438 VDD B12 INVB12 B13 INVB13 PCEN ICV_5 $T=-1695 -1270 0 0 $X=-2605 $Y=-1700
X439 VDD B14 INVB14 B15 INVB15 PCEN ICV_5 $T=7225 -1270 0 0 $X=6315 $Y=-1700
X440 VDD 361 O1 337 O0 GND 370 346 ICV_8 $T=-55075 -63750 1 180 $X=-56165 $Y=-64880
X441 VDD 409 O3 385 O2 GND 418 394 ICV_8 $T=-46155 -63750 1 180 $X=-47245 $Y=-64880
X442 VDD 457 O5 433 O4 GND 466 442 ICV_8 $T=-37235 -63750 1 180 $X=-38325 $Y=-64880
X443 VDD 505 O7 481 O6 GND 514 490 ICV_8 $T=-28315 -63750 1 180 $X=-29405 $Y=-64880
X444 VDD 553 O9 529 O8 GND 562 538 ICV_8 $T=-19395 -63750 1 180 $X=-20485 $Y=-64880
X445 VDD 601 O11 577 O10 GND 610 586 ICV_8 $T=-10475 -63750 1 180 $X=-11565 $Y=-64880
X446 VDD 649 O13 625 O12 GND 658 634 ICV_8 $T=-1555 -63750 1 180 $X=-2645 $Y=-64880
X447 VDD 697 O15 673 O14 GND 706 682 ICV_8 $T=7365 -63750 1 180 $X=6275 $Y=-64880
X448 GND VDD 327 338 351 362 375 386 399 410 423 434 447 458 471 482 495 506 519 530
+ 543 554 567 578 591 602 615 626 639 650 663 674 687 698
+ ICV_15 $T=-55255 -49230 0 0 $X=-56775 $Y=-49580
X449 GND VDD 328 339 352 363 376 387 400 411 424 435 448 459 472 483 496 507 520 531
+ 544 555 568 579 592 603 616 627 640 651 664 675 688 699
+ ICV_15 $T=-55255 -43190 0 0 $X=-56775 $Y=-43540
X450 GND VDD 329 340 353 364 377 388 401 412 425 436 449 460 473 484 497 508 521 532
+ 545 556 569 580 593 604 617 628 641 652 665 676 689 700
+ ICV_15 $T=-55255 -37150 0 0 $X=-56775 $Y=-37500
X451 GND VDD 330 341 354 365 378 389 402 413 426 437 450 461 474 485 498 509 522 533
+ 546 557 570 581 594 605 618 629 642 653 666 677 690 701
+ ICV_15 $T=-55255 -31110 0 0 $X=-56775 $Y=-31460
X452 GND VDD 331 342 355 366 379 390 403 414 427 438 451 462 475 486 499 510 523 534
+ 547 558 571 582 595 606 619 630 643 654 667 678 691 702
+ ICV_15 $T=-55255 -25070 0 0 $X=-56775 $Y=-25420
X453 GND VDD 332 343 356 367 380 391 404 415 428 439 452 463 476 487 500 511 524 535
+ 548 559 572 583 596 607 620 631 644 655 668 679 692 703
+ ICV_15 $T=-55255 -19030 0 0 $X=-56775 $Y=-19380
X454 GND VDD 333 344 357 368 381 392 405 416 429 440 453 464 477 488 501 512 525 536
+ 549 560 573 584 597 608 621 632 645 656 669 680 693 704
+ ICV_15 $T=-55255 -12990 0 0 $X=-56775 $Y=-13340
X455 GND VDD 334 345 358 369 382 393 406 417 430 441 454 465 478 489 502 513 526 537
+ 550 561 574 585 598 609 622 633 646 657 670 681 694 705
+ ICV_15 $T=-55255 -6950 0 0 $X=-56775 $Y=-7300
X456 GND 310 309 n18_CDNS_6737959159723 $T=-60915 -75550 0 0 $X=-61575 $Y=-76680
X457 GND CLKREG 310 n18_CDNS_6737959159723 $T=-58975 -75550 0 0 $X=-59635 $Y=-76680
X458 VDD 310 309 p18_CDNS_6737959159726 $T=-60915 -72930 0 0 $X=-61825 $Y=-73360
X459 VDD CLKREG 310 p18_CDNS_6737959159726 $T=-58975 -72930 0 0 $X=-59885 $Y=-73360
X460 GND 24 58 MODE n18_CDNS_6737959159725 $T=-66235 -61790 1 0 $X=-66895 $Y=-62580
X461 GND ADD7 69 MODE n18_CDNS_6737959159725 $T=-62355 -60310 0 0 $X=-63015 $Y=-61440
X462 GND ADD6 70 MODE n18_CDNS_6737959159725 $T=-62355 -46550 1 0 $X=-63015 $Y=-47340
X463 GND ADD5 71 MODE n18_CDNS_6737959159725 $T=-62355 -45070 0 0 $X=-63015 $Y=-46200
X464 GND ADD4 72 MODE n18_CDNS_6737959159725 $T=-62355 -31310 1 0 $X=-63015 $Y=-32100
X465 GND ADD3 73 MODE n18_CDNS_6737959159725 $T=-62355 -29830 0 0 $X=-63015 $Y=-30960
X466 GND ADD2 74 MODE n18_CDNS_6737959159725 $T=-62355 -16070 1 0 $X=-63015 $Y=-16860
X467 GND ADD1 75 MODE n18_CDNS_6737959159725 $T=-62355 -14590 0 0 $X=-63015 $Y=-15720
X468 GND ADD0 76 MODE n18_CDNS_6737959159725 $T=-62355 -830 1 0 $X=-63015 $Y=-1620
X469 GND GND 69 50 n18_CDNS_6737959159725 $T=-59695 -60310 0 0 $X=-60355 $Y=-61440
X470 GND GND 70 51 n18_CDNS_6737959159725 $T=-59695 -46550 1 0 $X=-60355 $Y=-47340
X471 GND GND 71 52 n18_CDNS_6737959159725 $T=-59695 -45070 0 0 $X=-60355 $Y=-46200
X472 GND GND 72 53 n18_CDNS_6737959159725 $T=-59695 -31310 1 0 $X=-60355 $Y=-32100
X473 GND GND 73 54 n18_CDNS_6737959159725 $T=-59695 -29830 0 0 $X=-60355 $Y=-30960
X474 GND GND 74 55 n18_CDNS_6737959159725 $T=-59695 -16070 1 0 $X=-60355 $Y=-16860
X475 GND GND 75 56 n18_CDNS_6737959159725 $T=-59695 -14590 0 0 $X=-60355 $Y=-15720
X476 GND 311 24 n18_CDNS_673795915970 $T=-60915 -61790 1 0 $X=-61575 $Y=-63020
X477 GND 186 196 185 ICV_16 $T=-96335 650 0 0 $X=-96995 $Y=-480
X478 GND 239 250 229 ICV_16 $T=-83595 -60310 0 0 $X=-84255 $Y=-61440
X479 GND 34 249 238 ICV_16 $T=-82755 650 0 0 $X=-83415 $Y=-480
X480 GND 289 306 279 ICV_16 $T=-71455 -75550 0 0 $X=-72115 $Y=-76680
X481 GND 312 PCEN 25 ICV_16 $T=-60915 650 0 0 $X=-61575 $Y=-480
X482 VDD 306 289 p18_CDNS_6737959159719 $T=-69515 -71170 0 0 $X=-70425 $Y=-71600
X483 VDD 249 267 34 ICV_17 $T=-80815 5030 0 0 $X=-81725 $Y=4600
X484 VDD 311 SAEN 24 ICV_17 $T=-60915 -66170 1 0 $X=-61825 $Y=-69060
X485 VDD 312 PCEN 25 ICV_17 $T=-60915 5030 0 0 $X=-61825 $Y=4600
X486 VDD MODE 735 p18_CDNS_6737959159720 $T=-66235 -67050 1 0 $X=-67145 $Y=-69060
X487 VDD 25 MODE 37 ICV_18 $T=-66235 5910 0 0 $X=-67145 $Y=5480
X488 VDD ADD7 MODE 40 ICV_18 $T=-62355 -55050 0 0 $X=-63265 $Y=-55480
X489 VDD ADD6 MODE 41 ICV_18 $T=-62355 -51810 1 0 $X=-63265 $Y=-53820
X490 VDD ADD5 MODE 42 ICV_18 $T=-62355 -39810 0 0 $X=-63265 $Y=-40240
X491 VDD ADD4 MODE 43 ICV_18 $T=-62355 -36570 1 0 $X=-63265 $Y=-38580
X492 VDD ADD3 MODE 44 ICV_18 $T=-62355 -24570 0 0 $X=-63265 $Y=-25000
X493 VDD ADD2 MODE 45 ICV_18 $T=-62355 -21330 1 0 $X=-63265 $Y=-23340
X494 VDD ADD1 MODE 46 ICV_18 $T=-62355 -9330 0 0 $X=-63265 $Y=-9760
X495 VDD ADD0 MODE 47 ICV_18 $T=-62355 -6090 1 0 $X=-63265 $Y=-8100
X496 GND 187 25 n18_CDNS_6737959159717 $T=-95355 -60210 0 0 $X=-96055 $Y=-61440
X497 GND 26 187 n18_CDNS_6737959159717 $T=-93335 -60210 0 0 $X=-94035 $Y=-61440
X498 GND 258 250 n18_CDNS_6737959159717 $T=-79675 -60210 0 0 $X=-80375 $Y=-61440
X499 GND 265 257 n18_CDNS_6737959159717 $T=-79675 -930 1 0 $X=-80375 $Y=-1500
X500 GND 278 267 n18_CDNS_6737959159717 $T=-76895 750 0 0 $X=-77595 $Y=-480
X501 GND 280 269 n18_CDNS_6737959159717 $T=-75035 -60210 0 0 $X=-75735 $Y=-61440
X502 GND 287 276 n18_CDNS_6737959159717 $T=-75035 -930 1 0 $X=-75735 $Y=-1500
X503 GND 36 34 n18_CDNS_6737959159717 $T=-72255 -61890 1 0 $X=-72955 $Y=-62460
X504 GND 37 288 n18_CDNS_6737959159717 $T=-72255 750 0 0 $X=-72955 $Y=-480
X505 GND 38 GND n18_CDNS_6737959159717 $T=-70235 -61890 1 0 $X=-70935 $Y=-62460
X506 GND 39 VDD n18_CDNS_6737959159717 $T=-70235 750 0 0 $X=-70935 $Y=-480
X507 GND 48 MODE n18_CDNS_6737959159717 $T=-68215 -61890 1 0 $X=-68915 $Y=-62460
X508 GND 49 MODE n18_CDNS_6737959159717 $T=-68215 750 0 0 $X=-68915 $Y=-480
X509 GND 307 306 n18_CDNS_6737959159717 $T=-67535 -75450 0 0 $X=-68235 $Y=-76680
X510 GND 57 2 n18_CDNS_6737959159717 $T=-66355 -930 1 0 $X=-67055 $Y=-1500
X511 GND 61 MODE n18_CDNS_6737959159717 $T=-64335 -60210 0 0 $X=-65035 $Y=-61440
X512 GND 68 MODE n18_CDNS_6737959159717 $T=-64335 -930 1 0 $X=-65035 $Y=-1500
X513 GND 309 308 n18_CDNS_6737959159717 $T=-62895 -75450 0 0 $X=-63595 $Y=-76680
X514 GND 269 26 712 n18_CDNS_6737959159722 $T=-77265 -60310 0 0 $X=-77585 $Y=-61440
X515 GND 270 27 713 n18_CDNS_6737959159722 $T=-77265 -46550 1 0 $X=-77585 $Y=-47340
X516 GND 271 28 714 n18_CDNS_6737959159722 $T=-77265 -45070 0 0 $X=-77585 $Y=-46200
X517 GND 272 29 715 n18_CDNS_6737959159722 $T=-77265 -31310 1 0 $X=-77585 $Y=-32100
X518 GND 273 30 716 n18_CDNS_6737959159722 $T=-77265 -29830 0 0 $X=-77585 $Y=-30960
X519 GND 274 31 717 n18_CDNS_6737959159722 $T=-77265 -16070 1 0 $X=-77585 $Y=-16860
X520 GND 275 32 718 n18_CDNS_6737959159722 $T=-77265 -14590 0 0 $X=-77585 $Y=-15720
X521 GND 291 281 719 n18_CDNS_6737959159722 $T=-72625 -46550 1 0 $X=-72945 $Y=-47340
X522 GND 292 282 720 n18_CDNS_6737959159722 $T=-72625 -45070 0 0 $X=-72945 $Y=-46200
X523 GND 293 283 721 n18_CDNS_6737959159722 $T=-72625 -31310 1 0 $X=-72945 $Y=-32100
X524 GND 294 284 722 n18_CDNS_6737959159722 $T=-72625 -29830 0 0 $X=-72945 $Y=-30960
X525 GND 295 285 723 n18_CDNS_6737959159722 $T=-72625 -16070 1 0 $X=-72945 $Y=-16860
X526 GND 296 286 724 n18_CDNS_6737959159722 $T=-72625 -14590 0 0 $X=-72945 $Y=-15720
X527 GND 308 307 725 n18_CDNS_6737959159722 $T=-65125 -75550 0 0 $X=-65445 $Y=-76680
X528 GND 258 712 n18_CDNS_6737959159724 $T=-77695 -60310 0 0 $X=-78355 $Y=-61440
X529 GND 259 713 n18_CDNS_6737959159724 $T=-77695 -46550 1 0 $X=-78355 $Y=-47340
X530 GND 260 714 n18_CDNS_6737959159724 $T=-77695 -45070 0 0 $X=-78355 $Y=-46200
X531 GND 261 715 n18_CDNS_6737959159724 $T=-77695 -31310 1 0 $X=-78355 $Y=-32100
X532 GND 262 716 n18_CDNS_6737959159724 $T=-77695 -29830 0 0 $X=-78355 $Y=-30960
X533 GND 263 717 n18_CDNS_6737959159724 $T=-77695 -16070 1 0 $X=-78355 $Y=-16860
X534 GND 264 718 n18_CDNS_6737959159724 $T=-77695 -14590 0 0 $X=-78355 $Y=-15720
X535 GND 265 708 n18_CDNS_6737959159724 $T=-77695 -830 1 0 $X=-78355 $Y=-1620
X536 GND 1 710 n18_CDNS_6737959159724 $T=-73055 -60310 0 0 $X=-73715 $Y=-61440
X537 GND 6 719 n18_CDNS_6737959159724 $T=-73055 -46550 1 0 $X=-73715 $Y=-47340
X538 GND 5 720 n18_CDNS_6737959159724 $T=-73055 -45070 0 0 $X=-73715 $Y=-46200
X539 GND 7 721 n18_CDNS_6737959159724 $T=-73055 -31310 1 0 $X=-73715 $Y=-32100
X540 GND 8 722 n18_CDNS_6737959159724 $T=-73055 -29830 0 0 $X=-73715 $Y=-30960
X541 GND 4 723 n18_CDNS_6737959159724 $T=-73055 -16070 1 0 $X=-73715 $Y=-16860
X542 GND 3 724 n18_CDNS_6737959159724 $T=-73055 -14590 0 0 $X=-73715 $Y=-15720
X543 GND 2 711 n18_CDNS_6737959159724 $T=-73055 -830 1 0 $X=-73715 $Y=-1620
X544 GND 60 725 n18_CDNS_6737959159724 $T=-65555 -75550 0 0 $X=-66215 $Y=-76680
X545 VDD 176 CLK p18_CDNS_6737959159718 $T=-103085 -48080 1 270 $X=-105095 $Y=-49170
X546 VDD 177 CLK p18_CDNS_6737959159718 $T=-103085 -43440 1 270 $X=-105095 $Y=-44530
X547 VDD 178 CLK p18_CDNS_6737959159718 $T=-103085 -38800 1 270 $X=-105095 $Y=-39890
X548 VDD 179 CLK p18_CDNS_6737959159718 $T=-103085 -34160 1 270 $X=-105095 $Y=-35250
X549 VDD 180 CLK p18_CDNS_6737959159718 $T=-103085 -29520 1 270 $X=-105095 $Y=-30610
X550 VDD 181 CLK p18_CDNS_6737959159718 $T=-103085 -24880 1 270 $X=-105095 $Y=-25970
X551 VDD 288 CLK p18_CDNS_6737959159718 $T=-74915 5910 0 0 $X=-75825 $Y=5480
X552 VDD 308 60 p18_CDNS_6737959159718 $T=-65555 -70290 0 0 $X=-66465 $Y=-70720
X553 GND 260 259 252 251 ICV_19 $T=-79675 -46650 1 0 $X=-80375 $Y=-47220
X554 GND 262 261 254 253 ICV_19 $T=-79675 -31410 1 0 $X=-80375 $Y=-31980
X555 GND 264 263 256 255 ICV_19 $T=-79675 -16170 1 0 $X=-80375 $Y=-16740
X556 GND 282 281 271 270 ICV_19 $T=-75035 -46650 1 0 $X=-75735 $Y=-47220
X557 GND 284 283 273 272 ICV_19 $T=-75035 -31410 1 0 $X=-75735 $Y=-31980
X558 GND 286 285 275 274 ICV_19 $T=-75035 -16170 1 0 $X=-75735 $Y=-16740
X559 GND 189 188 28 27 25 25 189 188 ICV_20 $T=-95355 -46650 1 0 $X=-96055 $Y=-47220
X560 GND 191 190 30 29 25 25 191 190 ICV_20 $T=-95355 -31410 1 0 $X=-96055 $Y=-31980
X561 GND 193 192 32 31 25 25 193 192 ICV_20 $T=-95355 -16170 1 0 $X=-96055 $Y=-16740
X562 GND 300 299 42 41 292 291 300 299 ICV_20 $T=-70395 -46650 1 0 $X=-71095 $Y=-47220
X563 GND 302 301 44 43 294 293 302 301 ICV_20 $T=-70395 -31410 1 0 $X=-71095 $Y=-31980
X564 GND 304 303 46 45 296 295 304 303 ICV_20 $T=-70395 -16170 1 0 $X=-71095 $Y=-16740
X565 GND 52 51 63 62 5 6 MODE MODE ICV_20 $T=-66355 -46650 1 0 $X=-67055 $Y=-47220
X566 GND 54 53 65 64 8 7 MODE MODE ICV_20 $T=-66355 -31410 1 0 $X=-67055 $Y=-31980
X567 GND 56 55 67 66 3 4 MODE MODE ICV_20 $T=-66355 -16170 1 0 $X=-67055 $Y=-16740
X568 VDD 258 259 250 251 ICV_21 $T=-79675 -54610 0 0 $X=-80585 $Y=-55040
X569 VDD 260 261 252 253 ICV_21 $T=-79675 -39370 0 0 $X=-80585 $Y=-39800
X570 VDD 262 263 254 255 ICV_21 $T=-79675 -24130 0 0 $X=-80585 $Y=-24560
X571 VDD 264 265 256 257 ICV_21 $T=-79675 -8890 0 0 $X=-80585 $Y=-9320
X572 VDD 280 281 269 270 ICV_21 $T=-75035 -54610 0 0 $X=-75945 $Y=-55040
X573 VDD 282 283 271 272 ICV_21 $T=-75035 -39370 0 0 $X=-75945 $Y=-39800
X574 VDD 284 285 273 274 ICV_21 $T=-75035 -24130 0 0 $X=-75945 $Y=-24560
X575 VDD 286 287 275 276 ICV_21 $T=-75035 -8890 0 0 $X=-75945 $Y=-9320
X576 VDD 187 188 26 27 25 25 187 188 ICV_22 $T=-95355 -54610 0 0 $X=-96265 $Y=-55040
X577 VDD 189 190 28 29 25 25 189 190 ICV_22 $T=-95355 -39370 0 0 $X=-96265 $Y=-39800
X578 VDD 191 192 30 31 25 25 191 192 ICV_22 $T=-95355 -24130 0 0 $X=-96265 $Y=-24560
X579 VDD 193 194 32 33 25 25 193 194 ICV_22 $T=-95355 -8890 0 0 $X=-96265 $Y=-9320
X580 VDD 298 299 40 41 290 291 298 299 ICV_22 $T=-70395 -54610 0 0 $X=-71305 $Y=-55040
X581 VDD 300 301 42 43 292 293 300 301 ICV_22 $T=-70395 -39370 0 0 $X=-71305 $Y=-39800
X582 VDD 302 303 44 45 294 295 302 303 ICV_22 $T=-70395 -24130 0 0 $X=-71305 $Y=-24560
X583 VDD 304 305 46 47 296 297 304 305 ICV_22 $T=-70395 -8890 0 0 $X=-71305 $Y=-9320
X584 VDD 50 51 61 62 1 6 MODE MODE ICV_22 $T=-66355 -54610 0 0 $X=-67265 $Y=-55040
X585 VDD 52 53 63 64 5 7 MODE MODE ICV_22 $T=-66355 -39370 0 0 $X=-67265 $Y=-39800
X586 VDD 54 55 65 66 8 4 MODE MODE ICV_22 $T=-66355 -24130 0 0 $X=-67265 $Y=-24560
X587 VDD 56 57 67 68 3 2 MODE MODE ICV_22 $T=-66355 -8890 0 0 $X=-67265 $Y=-9320
X588 VDD 269 270 258 259 ICV_23 $T=-77695 -55050 0 0 $X=-78605 $Y=-55480
X589 VDD 271 272 260 261 ICV_23 $T=-77695 -39810 0 0 $X=-78605 $Y=-40240
X590 VDD 273 274 262 263 ICV_23 $T=-77695 -24570 0 0 $X=-78605 $Y=-25000
X591 VDD 275 276 264 265 ICV_23 $T=-77695 -9330 0 0 $X=-78605 $Y=-9760
X592 VDD 290 291 1 6 ICV_23 $T=-73055 -55050 0 0 $X=-73965 $Y=-55480
X593 VDD 292 293 5 7 ICV_23 $T=-73055 -39810 0 0 $X=-73965 $Y=-40240
X594 VDD 294 295 8 4 ICV_23 $T=-73055 -24570 0 0 $X=-73965 $Y=-25000
X595 VDD 296 297 3 2 ICV_23 $T=-73055 -9330 0 0 $X=-73965 $Y=-9760
X596 GND 201 200 211 210 28 27 ICV_25 $T=-91355 -46550 1 0 $X=-92015 $Y=-47780
X597 GND 203 202 213 212 30 29 ICV_25 $T=-91355 -31310 1 0 $X=-92015 $Y=-32540
X598 GND 205 204 215 214 32 31 ICV_25 $T=-91355 -16070 1 0 $X=-92015 $Y=-17300
X599 GND 221 220 231 230 211 210 ICV_25 $T=-87475 -46550 1 0 $X=-88135 $Y=-47780
X600 GND 223 222 233 232 213 212 ICV_25 $T=-87475 -31310 1 0 $X=-88135 $Y=-32540
X601 GND 225 224 235 234 215 214 ICV_25 $T=-87475 -16070 1 0 $X=-88135 $Y=-17300
X602 GND 241 240 252 251 231 230 ICV_25 $T=-83595 -46550 1 0 $X=-84255 $Y=-47780
X603 GND 243 242 254 253 233 232 ICV_25 $T=-83595 -31310 1 0 $X=-84255 $Y=-32540
X604 GND 245 244 256 255 235 234 ICV_25 $T=-83595 -16070 1 0 $X=-84255 $Y=-17300
X605 VDD 239 250 240 251 229 230 ICV_26 $T=-83595 -55930 0 0 $X=-84505 $Y=-56360
X606 VDD 241 252 242 253 231 232 ICV_26 $T=-83595 -40690 0 0 $X=-84505 $Y=-41120
X607 VDD 243 254 244 255 233 234 ICV_26 $T=-83595 -25450 0 0 $X=-84505 $Y=-25880
X608 VDD 245 256 246 257 235 236 ICV_26 $T=-83595 -10210 0 0 $X=-84505 $Y=-10640
X609 GND 199 209 219 229 26 ICV_27 $T=-91355 -60310 0 0 $X=-92015 $Y=-61440
X610 GND 208 218 228 238 198 ICV_27 $T=-90515 650 0 0 $X=-91175 $Y=-480
X611 GND 143 144 145 146 147 148 149 150 24 ICV_28 $T=-149055 -75550 0 0 $X=-149715 $Y=-76680
X612 GND 151 152 153 154 155 156 157 158 150 ICV_28 $T=-133535 -75550 0 0 $X=-134195 $Y=-76680
X613 GND 159 160 161 162 164 166 168 170 158 ICV_28 $T=-118015 -75550 0 0 $X=-118675 $Y=-76680
X614 GND 163 165 167 169 171 173 175 185 CLK ICV_28 $T=-111855 650 0 0 $X=-112515 $Y=-480
X615 GND 172 174 184 60 195 197 207 217 170 ICV_28 $T=-102495 -75550 0 0 $X=-103155 $Y=-76680
X616 GND 227 237 247 248 266 268 277 279 217 ICV_28 $T=-86975 -75550 0 0 $X=-87635 $Y=-76680
X617 VDD 143 144 145 146 147 148 149 150 24 ICV_30 $T=-149055 -71170 0 0 $X=-149965 $Y=-71600
X618 VDD 151 152 153 154 155 156 157 158 150 ICV_30 $T=-133535 -71170 0 0 $X=-134445 $Y=-71600
X619 VDD 159 160 161 162 164 166 168 170 158 ICV_30 $T=-118015 -71170 0 0 $X=-118925 $Y=-71600
X620 VDD 163 165 167 169 171 173 175 185 CLK ICV_30 $T=-111855 5030 0 0 $X=-112765 $Y=4600
X621 VDD 172 174 184 60 195 197 207 217 170 ICV_30 $T=-102495 -71170 0 0 $X=-103405 $Y=-71600
X622 VDD 186 196 198 208 218 228 238 34 185 ICV_30 $T=-96335 5030 0 0 $X=-97245 $Y=4600
X623 VDD 227 237 247 248 266 268 277 279 217 ICV_30 $T=-86975 -71170 0 0 $X=-87885 $Y=-71600
X624 VDD 199 200 209 210 219 220 229 230 26 27 ICV_31 $T=-91355 -55930 0 0 $X=-92265 $Y=-56360
X625 VDD 201 202 211 212 221 222 231 232 28 29 ICV_31 $T=-91355 -40690 0 0 $X=-92265 $Y=-41120
X626 VDD 203 204 213 214 223 224 233 234 30 31 ICV_31 $T=-91355 -25450 0 0 $X=-92265 $Y=-25880
X627 VDD 205 206 215 216 225 226 235 236 32 33 ICV_31 $T=-91355 -10210 0 0 $X=-92265 $Y=-10640
X628 GND 1 176 15 CLK ICV_32 $T=-97925 -50740 1 270 $X=-98615 $Y=-51620
X629 GND 6 177 18 CLK ICV_32 $T=-97925 -46100 1 270 $X=-98615 $Y=-46980
X630 GND 5 178 19 CLK ICV_32 $T=-97925 -41460 1 270 $X=-98615 $Y=-42340
X631 GND 7 179 20 CLK ICV_32 $T=-97925 -36820 1 270 $X=-98615 $Y=-37700
X632 GND 8 180 21 CLK ICV_32 $T=-97925 -32180 1 270 $X=-98615 $Y=-33060
X633 GND 4 181 22 CLK ICV_32 $T=-97925 -27540 1 270 $X=-98615 $Y=-28420
X634 GND 3 182 16 CLK ICV_32 $T=-97925 -22900 1 270 $X=-98615 $Y=-23780
X635 GND 2 183 17 CLK ICV_32 $T=-97925 -18260 1 270 $X=-98615 $Y=-19140
X636 VDD 13 746 p18_CDNS_673795915971 $T=-106765 -26460 0 270 $X=-107195 $Y=-27195
X637 VDD A0 747 p18_CDNS_673795915971 $T=-106765 -22840 0 270 $X=-107195 $Y=-23575
X638 VDD 13 734 p18_CDNS_673795915971 $T=-106765 -19220 0 270 $X=-107195 $Y=-19955
X639 VDD A0 748 p18_CDNS_673795915971 $T=-106765 -15600 0 270 $X=-107195 $Y=-16335
X640 VDD 14 727 726 p18_CDNS_6737959159729 $T=-106765 -41370 0 270 $X=-107195 $Y=-42105
X641 VDD A1 732 749 p18_CDNS_6737959159729 $T=-106765 -30510 0 270 $X=-107195 $Y=-31245
X642 VDD 14 746 750 p18_CDNS_6737959159729 $T=-106765 -26890 0 270 $X=-107195 $Y=-27625
X643 VDD 14 747 751 p18_CDNS_6737959159729 $T=-106765 -23270 0 270 $X=-107195 $Y=-24005
X644 VDD A1 748 752 p18_CDNS_6737959159729 $T=-106765 -16030 0 270 $X=-107195 $Y=-16765
X645 VDD 20 12 749 p18_CDNS_6737959159728 $T=-106765 -30940 0 270 $X=-107195 $Y=-32030
X646 VDD 21 A2 750 p18_CDNS_6737959159728 $T=-106765 -27320 0 270 $X=-107195 $Y=-28410
X647 VDD 22 A2 751 p18_CDNS_6737959159728 $T=-106765 -23700 0 270 $X=-107195 $Y=-24790
X648 VDD 16 A2 733 p18_CDNS_6737959159728 $T=-106765 -20080 0 270 $X=-107195 $Y=-21170
X649 VDD 17 A2 752 p18_CDNS_6737959159728 $T=-106765 -16460 0 270 $X=-107195 $Y=-17550
X650 GND GND 12 A2 n18_CDNS_6737959159727 $T=-110435 -42540 1 270 $X=-111005 $Y=-43420
X651 GND GND 14 A1 n18_CDNS_6737959159727 $T=-110435 -40520 1 270 $X=-111005 $Y=-41400
X652 GND 15 GND 12 n18_CDNS_6737959159727 $T=-108935 -42540 0 270 $X=-110075 $Y=-43420
X653 GND 18 GND A0 n18_CDNS_6737959159727 $T=-108935 -37320 0 270 $X=-110075 $Y=-38200
X654 GND 19 GND 12 n18_CDNS_6737959159727 $T=-108935 -35300 0 270 $X=-110075 $Y=-36180
X655 GND 19 GND 13 n18_CDNS_6737959159727 $T=-108935 -33700 0 270 $X=-110075 $Y=-34580
X656 GND 20 GND 12 n18_CDNS_6737959159727 $T=-108935 -31680 0 270 $X=-110075 $Y=-32560
X657 GND 20 GND A0 n18_CDNS_6737959159727 $T=-108935 -30080 0 270 $X=-110075 $Y=-30960
X658 GND 21 GND A2 n18_CDNS_6737959159727 $T=-108935 -28060 0 270 $X=-110075 $Y=-28940
X659 GND 21 GND 13 n18_CDNS_6737959159727 $T=-108935 -26460 0 270 $X=-110075 $Y=-27340
X660 GND 22 GND A2 n18_CDNS_6737959159727 $T=-108935 -24440 0 270 $X=-110075 $Y=-25320
X661 GND 22 GND A0 n18_CDNS_6737959159727 $T=-108935 -22840 0 270 $X=-110075 $Y=-23720
X662 GND 16 GND A2 n18_CDNS_6737959159727 $T=-108935 -20820 0 270 $X=-110075 $Y=-21700
X663 GND 16 GND 13 n18_CDNS_6737959159727 $T=-108935 -19220 0 270 $X=-110075 $Y=-20100
X664 GND 17 GND A2 n18_CDNS_6737959159727 $T=-108935 -17200 0 270 $X=-110075 $Y=-18080
X665 GND 17 GND A0 n18_CDNS_6737959159727 $T=-108935 -15600 0 270 $X=-110075 $Y=-16480
.ENDS
***************************************

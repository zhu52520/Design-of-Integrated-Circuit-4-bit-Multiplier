* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_672414149280 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_672414149281 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672414149283 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672414149284 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 4 3 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672414149282 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT CSA_B INVCOUT COUT B A S INVCI CI GND VDD
** N=23 EP=9 IP=77 FDC=40
M0 6 CI INVCOUT GND NM L=1.8e-07 W=4.4e-07 $X=4005 $Y=-22185 $D=0
M1 11 CI COUT GND NM L=1.8e-07 W=4.4e-07 $X=5945 $Y=-22185 $D=0
M2 GND 6 11 GND NM L=1.8e-07 W=4.4e-07 $X=6665 $Y=-22185 $D=0
M3 GND 7 10 GND NM L=1.8e-07 W=4.4e-07 $X=6865 $Y=-18485 $D=0
M4 6 A GND GND NM L=1.8e-07 W=2.2e-07 $X=7425 $Y=-22085 $D=0
M5 20 B GND GND NM L=1.8e-07 W=4.4e-07 $X=7585 $Y=-18485 $D=0
M6 7 A 20 GND NM L=1.8e-07 W=4.4e-07 $X=8015 $Y=-18485 $D=0
M7 GND B 6 GND NM L=1.8e-07 W=2.2e-07 $X=8225 $Y=-22085 $D=0
M8 14 7 12 GND NM L=1.8e-07 W=4.4e-07 $X=9955 $Y=-18485 $D=0
M9 21 A 15 GND NM L=1.8e-07 W=4.4e-07 $X=10205 $Y=-22185 $D=0
M10 GND B 21 GND NM L=1.8e-07 W=4.4e-07 $X=10635 $Y=-22185 $D=0
M11 GND B 14 GND NM L=1.8e-07 W=4.4e-07 $X=10675 $Y=-18485 $D=0
M12 15 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=11395 $Y=-22085 $D=0
M13 14 A GND GND NM L=1.8e-07 W=4.4e-07 $X=11395 $Y=-18485 $D=0
M14 18 15 GND GND NM L=1.8e-07 W=4.4e-07 $X=13375 $Y=-22185 $D=0
M15 19 12 GND GND NM L=1.8e-07 W=4.4e-07 $X=13375 $Y=-18485 $D=0
M16 S CI 18 GND NM L=1.8e-07 W=4.4e-07 $X=14135 $Y=-22185 $D=0
M17 10 CI COUT VDD PM L=1.8e-07 W=4.4e-07 $X=6065 $Y=-15040 $D=4
M18 VDD 6 11 VDD PM L=1.8e-07 W=8.8e-07 $X=6865 $Y=-25630 $D=4
M19 7 B VDD VDD PM L=1.8e-07 W=4.4e-07 $X=7585 $Y=-15040 $D=4
M20 12 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=10245 $Y=-15040 $D=4
M21 13 B VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10675 $Y=-25630 $D=4
M22 S INVCI 18 VDD PM L=1.8e-07 W=4.4e-07 $X=14095 $Y=-25630 $D=4
M23 S CI 19 VDD PM L=1.8e-07 W=4.4e-07 $X=14135 $Y=-15040 $D=4
X24 GND 7 INVCOUT INVCI n18_CDNS_672414149280 $T=4295 -18485 1 180 $X=3455 $Y=-20505
X25 GND 10 COUT INVCI n18_CDNS_672414149280 $T=6245 -18485 1 180 $X=5405 $Y=-20505
X26 GND S 19 INVCI n18_CDNS_672414149280 $T=14315 -18485 1 180 $X=13475 $Y=-20505
X27 VDD 10 VDD 7 p18_CDNS_672414149281 $T=6825 -15480 0 0 $X=5915 $Y=-15910
X28 VDD 13 VDD A p18_CDNS_672414149281 $T=9955 -24750 1 0 $X=9045 $Y=-26980
X29 VDD 13 15 6 p18_CDNS_672414149281 $T=11395 -24750 1 0 $X=10485 $Y=-26980
X30 VDD VDD 18 15 p18_CDNS_672414149281 $T=13335 -24750 1 0 $X=12425 $Y=-26980
X31 VDD VDD 19 12 p18_CDNS_672414149281 $T=13375 -15480 0 0 $X=12465 $Y=-15910
X32 VDD 6 B 22 p18_CDNS_672414149283 $T=8015 -24750 1 0 $X=7460 $Y=-26980
X33 VDD VDD A 23 p18_CDNS_672414149283 $T=11435 -15480 0 0 $X=10880 $Y=-15910
X34 VDD VDD A 22 p18_CDNS_672414149284 $T=7585 -24750 1 0 $X=6675 $Y=-26980
X35 VDD 12 B 23 p18_CDNS_672414149284 $T=11005 -15480 0 0 $X=10095 $Y=-15910
X36 VDD INVCOUT 7 CI p18_CDNS_672414149282 $T=4115 -15040 0 0 $X=3205 $Y=-15470
X37 VDD 6 INVCOUT INVCI p18_CDNS_672414149282 $T=4345 -25190 0 180 $X=3255 $Y=-26980
X38 VDD 11 COUT INVCI p18_CDNS_672414149282 $T=6285 -25190 0 180 $X=5195 $Y=-26980
X39 VDD 7 VDD A p18_CDNS_672414149282 $T=8305 -15040 0 0 $X=7395 $Y=-15470
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_6738713766025 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766022 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 1 3 2 1 PM L=1.8e-07 W=3.3e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766029 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766021 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766023 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766018 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 5 6 n18_CDNS_6738713766023 $T=0 -1660 0 0 $X=-660 $Y=-2010
X1 3 4 5 6 n18_CDNS_6738713766018 $T=0 0 0 0 $X=-660 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766016 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766017 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=16 FDC=4
X0 1 2 1 6 n18_CDNS_6738713766016 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 1 3 7 n18_CDNS_6738713766016 $T=2020 0 0 0 $X=1360 $Y=-1130
X2 1 2 4 8 n18_CDNS_6738713766017 $T=0 2900 0 0 $X=-660 $Y=2550
X3 1 5 3 8 n18_CDNS_6738713766017 $T=2020 2900 0 0 $X=1360 $Y=2550
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=8
X0 1 2 5 3 4 10 12 11 ICV_2 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 9 7 8 13 14 11 ICV_2 $T=4460 0 0 0 $X=3800 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376605 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4
** N=5 EP=4 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_673871376605 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 1 4 p18_CDNS_673871376605 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6
** N=7 EP=6 IP=10 FDC=4
X0 1 2 3 6 ICV_4 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 6 ICV_4 $T=4460 0 0 0 $X=3550 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766020 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4
** N=5 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_6738713766020 $T=-2020 0 0 0 $X=-2930 $Y=-1130
X1 1 3 2 p18_CDNS_6738713766020 $T=0 0 0 0 $X=-910 $Y=-1130
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766024 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766019 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_6738713766024 $T=-2020 0 0 0 $X=-2720 $Y=-350
X1 1 3 2 n18_CDNS_6738713766019 $T=0 0 0 0 $X=-700 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=8
X0 1 2 3 7 ICV_6 $T=-4460 0 0 0 $X=-7390 $Y=-1130
X1 1 4 5 8 ICV_6 $T=0 0 0 0 $X=-2930 $Y=-1130
X2 6 2 3 7 ICV_7 $T=-4460 1650 0 0 $X=-7180 $Y=1300
X3 6 4 5 8 ICV_7 $T=0 1650 0 0 $X=-2720 $Y=1300
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766015 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766026 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 n18_CDNS_6738713766015 $T=0 0 0 0 $X=-1520 $Y=-350
X1 3 1 2 n18_CDNS_6738713766026 $T=2020 0 0 0 $X=1360 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_9 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 4 5 ICV_9 $T=4460 0 0 0 $X=2940 $Y=-350
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766028 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3
** N=3 EP=3 IP=8 FDC=2
X0 1 1 2 3 p18_CDNS_6738713766028 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 3 1 2 p18_CDNS_6738713766028 $T=2020 0 0 0 $X=1070 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_11 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 4 5 ICV_11 $T=4460 0 0 0 $X=3510 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=20 FDC=16
X0 1 2 3 4 5 ICV_10 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 6 7 8 9 ICV_10 $T=8920 0 0 0 $X=7400 $Y=-350
X2 10 2 3 4 5 ICV_12 $T=0 1950 0 0 $X=-950 $Y=1420
X3 10 6 7 8 9 ICV_12 $T=8920 1950 0 0 $X=7970 $Y=1420
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=20 FDC=32
X0 1 3 4 5 6 7 8 9 10 2 ICV_13 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 11 12 13 14 15 16 17 18 2 ICV_13 $T=17840 0 0 0 $X=16320 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=34 EP=34 IP=36 FDC=64
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_14 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 2 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_14 $T=35680 0 0 0 $X=34160 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766013 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766014 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=3.52e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766011 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673871376608 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673871376608 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 3 2 n18_CDNS_673871376608 $T=1940 0 0 0 $X=1280 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376609 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_673871376609 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 2 p18_CDNS_673871376609 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766010 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6738713766012 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4
** N=5 EP=4 IP=7 FDC=2
X0 1 3 5 p18_CDNS_6738713766010 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 2 4 5 p18_CDNS_6738713766012 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_673871376606 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673871376600 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673871376601 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376607 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673871376606 $T=0 -1680 1 0 $X=-700 $Y=-2250
X1 1 3 5 n18_CDNS_673871376606 $T=0 0 0 0 $X=-700 $Y=-1230
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_19 $T=0 0 0 0 $X=-700 $Y=-2250
X1 1 4 5 8 9 ICV_19 $T=2020 0 0 0 $X=1320 $Y=-2250
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_673871376605 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 1 3 5 p18_CDNS_673871376605 $T=0 2360 1 0 $X=-910 $Y=790
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_21 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 8 9 ICV_21 $T=2020 0 0 0 $X=1110 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 p18_CDNS_673871376607 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 p18_CDNS_673871376607 $T=0 3240 1 0 $X=-910 $Y=1230
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673871376608 $T=0 -1480 1 0 $X=-660 $Y=-2710
X1 1 3 5 n18_CDNS_673871376608 $T=0 0 0 0 $X=-660 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=4
X0 1 2 3 6 7 ICV_24 $T=0 0 0 0 $X=-660 $Y=-2710
X1 1 4 5 2 3 ICV_24 $T=1940 0 0 0 $X=1280 $Y=-2710
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7
** N=7 EP=7 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 7 ICV_17 $T=0 5000 1 0 $X=-910 $Y=2110
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_16 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 4 5 3 ICV_16 $T=3880 0 0 0 $X=3220 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=8
X0 1 2 3 4 5 10 ICV_27 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 7 8 9 5 ICV_27 $T=7760 0 0 0 $X=7100 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6
** N=7 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 3 ICV_17 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10
** N=11 EP=10 IP=14 FDC=8
X0 1 2 3 4 5 10 ICV_29 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 7 8 9 5 ICV_29 $T=7760 0 0 0 $X=6850 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=8
X0 1 2 4 3 5 10 11 ICV_26 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 8 7 9 4 5 ICV_26 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5
** N=6 EP=5 IP=10 FDC=3
X0 1 2 3 n18_CDNS_673871376606 $T=0 0 0 0 $X=-700 $Y=-1230
X1 1 3 4 6 n18_CDNS_673871376600 $T=-2230 -100 0 0 $X=-2550 $Y=-1230
X2 1 5 6 n18_CDNS_673871376601 $T=-2660 -100 0 0 $X=-3320 $Y=-1230
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376604 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376603 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 2 3 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673871376602 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6738713766027 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT SRAM_REG A2 A1 A0 GND CLK MODE CLKREG B0 INVB0 B1 INVB1 B2 INVB2 B3 INVB3 B4 INVB4 B5 INVB5 B6
+ INVB6 RST B7 INVB7 B8 INVB8 B9 INVB9 B10 INVB10 B11 INVB11 B12 INVB12 B13 INVB13 B14 INVB14 B15 INVB15
+ VDD ADD4 ADD3 SAEN ADD7 ADD6 ADD5 ADD2 ADD1 ADD0 PCEN D0 Q1 Q0 D1 Q3 Q2 D2 D3 Q5
+ Q4 D4 D5 Q7 Q6 D6 D7 Q9 Q8 D8 D9 Q11 Q10 D10 D11 Q13 Q12 D12 Q15 Q14
+ D13 D14 D15
** N=881 EP=83 IP=2653 FDC=1924
M0 GND A0 29 GND NM L=1.8e-07 W=2.2e-07 $X=-13265 $Y=2460 $D=0
M1 GND 30 31 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=-780 $D=0
M2 31 29 GND GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=20 $D=0
M3 34 28 GND GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=2040 $D=0
M4 GND 30 34 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=2840 $D=0
M5 GND A1 35 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=6460 $D=0
M6 GND A1 36 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=10080 $D=0
M7 GND 30 37 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=13700 $D=0
M8 GND 30 38 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=17320 $D=0
M9 GND A1 32 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=20940 $D=0
M10 GND A1 33 GND NM L=1.8e-07 W=2.2e-07 $X=-11545 $Y=24560 $D=0
M11 212 41 GND GND NM L=1.8e-07 W=2.2e-07 $X=2035 $Y=39990 $D=0
M12 49 212 GND GND NM L=1.8e-07 W=2.2e-07 $X=4055 $Y=39990 $D=0
M13 216 214 GND GND NM L=1.8e-07 W=8.8e-07 $X=4935 $Y=41790 $D=0
M14 224 49 GND GND NM L=1.8e-07 W=8.8e-07 $X=6035 $Y=39430 $D=0
M15 234 224 GND GND NM L=1.8e-07 W=8.8e-07 $X=7975 $Y=39430 $D=0
M16 244 234 GND GND NM L=1.8e-07 W=8.8e-07 $X=9915 $Y=39430 $D=0
M17 254 244 GND GND NM L=1.8e-07 W=8.8e-07 $X=11855 $Y=39430 $D=0
M18 264 254 GND GND NM L=1.8e-07 W=8.8e-07 $X=13795 $Y=39430 $D=0
M19 275 264 GND GND NM L=1.8e-07 W=8.8e-07 $X=15735 $Y=39430 $D=0
M20 285 267 GND GND NM L=1.8e-07 W=8.8e-07 $X=18515 $Y=41790 $D=0
M21 294 49 773 GND NM L=1.8e-07 W=4.4e-07 $X=20125 $Y=39870 $D=0
M22 774 CLK GND GND NM L=1.8e-07 W=4.4e-07 $X=22475 $Y=41790 $D=0
M23 306 296 774 GND NM L=1.8e-07 W=4.4e-07 $X=22905 $Y=41790 $D=0
M24 308 298 775 GND NM L=1.8e-07 W=4.4e-07 $X=24765 $Y=-19170 $D=0
M25 315 305 776 GND NM L=1.8e-07 W=4.4e-07 $X=24765 $Y=39870 $D=0
M26 316 308 GND GND NM L=1.8e-07 W=2.2e-07 $X=26995 $Y=-19070 $D=0
M27 323 315 GND GND NM L=1.8e-07 W=2.2e-07 $X=26995 $Y=39990 $D=0
M28 56 316 GND GND NM L=1.8e-07 W=2.2e-07 $X=29015 $Y=-19070 $D=0
M29 63 323 GND GND NM L=1.8e-07 W=2.2e-07 $X=29015 $Y=39990 $D=0
M30 66 1 GND GND NM L=1.8e-07 W=2.2e-07 $X=31035 $Y=-19070 $D=0
M31 75 MODE 41 GND NM L=1.8e-07 W=4.4e-07 $X=31155 $Y=41790 $D=0
M32 40 52 74 GND NM L=1.8e-07 W=4.4e-07 $X=31875 $Y=-21090 $D=0
M33 41 53 75 GND NM L=1.8e-07 W=4.4e-07 $X=31875 $Y=41790 $D=0
M34 74 54 GND GND NM L=1.8e-07 W=4.4e-07 $X=33815 $Y=-21090 $D=0
M35 75 55 GND GND NM L=1.8e-07 W=4.4e-07 $X=33815 $Y=41790 $D=0
M36 GND 64 74 GND NM L=1.8e-07 W=4.4e-07 $X=34535 $Y=-21090 $D=0
M37 GND 65 75 GND NM L=1.8e-07 W=4.4e-07 $X=34535 $Y=41790 $D=0
M38 ADD7 56 85 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=-19170 $D=0
M39 ADD6 57 86 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=-5850 $D=0
M40 ADD5 58 87 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=-3930 $D=0
M41 ADD4 59 88 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=9390 $D=0
M42 ADD3 60 89 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=11310 $D=0
M43 ADD2 61 90 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=24630 $D=0
M44 ADD1 62 91 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=26550 $D=0
M45 ADD0 63 92 GND NM L=1.8e-07 W=4.4e-07 $X=35755 $Y=39870 $D=0
M46 92 73 GND GND NM L=1.8e-07 W=4.4e-07 $X=37695 $Y=39870 $D=0
M47 SAEN 329 GND GND NM L=1.8e-07 W=8.8e-07 $X=38415 $Y=-21530 $D=0
M48 GND 77 85 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=-19170 $D=0
M49 GND 78 86 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=-5850 $D=0
M50 GND 79 87 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=-3930 $D=0
M51 GND 80 88 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=9390 $D=0
M52 GND 81 89 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=11310 $D=0
M53 GND 82 90 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=24630 $D=0
M54 GND 83 91 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=26550 $D=0
M55 GND 84 92 GND NM L=1.8e-07 W=4.4e-07 $X=38415 $Y=39870 $D=0
M56 777 365 GND GND NM L=1.8e-07 W=4.4e-07 $X=42135 $Y=-42825 $D=0
M57 778 366 GND GND NM L=1.8e-07 W=4.4e-07 $X=42135 $Y=-39125 $D=0
M58 Q1 CLKREG 777 GND NM L=1.8e-07 W=4.4e-07 $X=42565 $Y=-42825 $D=0
M59 Q0 CLKREG 778 GND NM L=1.8e-07 W=4.4e-07 $X=42565 $Y=-39125 $D=0
M60 GND D0 94 GND NM L=1.8e-07 W=2.2e-07 $X=42745 $Y=-26240 $D=0
M61 354 B0 342 GND NM L=1.8e-07 W=4.4e-07 $X=42785 $Y=-17660 $D=0
M62 98 94 GND GND NM L=1.8e-07 W=2.2e-07 $X=43545 $Y=-26240 $D=0
M63 779 CLKREG 365 GND NM L=1.8e-07 W=4.4e-07 $X=44505 $Y=-42825 $D=0
M64 780 CLKREG 366 GND NM L=1.8e-07 W=4.4e-07 $X=44505 $Y=-39125 $D=0
M65 GND 369 779 GND NM L=1.8e-07 W=4.4e-07 $X=44935 $Y=-42825 $D=0
M66 GND 370 780 GND NM L=1.8e-07 W=4.4e-07 $X=44935 $Y=-39125 $D=0
M67 369 382 GND GND NM L=1.8e-07 W=4.4e-07 $X=45655 $Y=-42825 $D=0
M68 370 383 GND GND NM L=1.8e-07 W=4.4e-07 $X=45655 $Y=-39125 $D=0
M69 GND RST 369 GND NM L=1.8e-07 W=4.4e-07 $X=46375 $Y=-42825 $D=0
M70 GND RST 370 GND NM L=1.8e-07 W=4.4e-07 $X=46375 $Y=-39125 $D=0
M71 GND D1 99 GND NM L=1.8e-07 W=2.2e-07 $X=47205 $Y=-26240 $D=0
M72 381 B1 371 GND NM L=1.8e-07 W=4.4e-07 $X=47245 $Y=-17660 $D=0
M73 102 99 GND GND NM L=1.8e-07 W=2.2e-07 $X=48005 $Y=-26240 $D=0
M74 GND 10 382 GND NM L=1.8e-07 W=2.2e-07 $X=48355 $Y=-42725 $D=0
M75 GND 9 383 GND NM L=1.8e-07 W=2.2e-07 $X=48355 $Y=-39005 $D=0
M76 781 409 GND GND NM L=1.8e-07 W=4.4e-07 $X=50335 $Y=-42825 $D=0
M77 782 410 GND GND NM L=1.8e-07 W=4.4e-07 $X=50335 $Y=-39125 $D=0
M78 Q3 CLKREG 781 GND NM L=1.8e-07 W=4.4e-07 $X=50765 $Y=-42825 $D=0
M79 Q2 CLKREG 782 GND NM L=1.8e-07 W=4.4e-07 $X=50765 $Y=-39125 $D=0
M80 GND D2 103 GND NM L=1.8e-07 W=2.2e-07 $X=51665 $Y=-26240 $D=0
M81 408 B2 398 GND NM L=1.8e-07 W=4.4e-07 $X=51705 $Y=-17660 $D=0
M82 106 103 GND GND NM L=1.8e-07 W=2.2e-07 $X=52465 $Y=-26240 $D=0
M83 783 CLKREG 409 GND NM L=1.8e-07 W=4.4e-07 $X=52705 $Y=-42825 $D=0
M84 784 CLKREG 410 GND NM L=1.8e-07 W=4.4e-07 $X=52705 $Y=-39125 $D=0
M85 GND 423 783 GND NM L=1.8e-07 W=4.4e-07 $X=53135 $Y=-42825 $D=0
M86 GND 424 784 GND NM L=1.8e-07 W=4.4e-07 $X=53135 $Y=-39125 $D=0
M87 423 434 GND GND NM L=1.8e-07 W=4.4e-07 $X=53855 $Y=-42825 $D=0
M88 424 435 GND GND NM L=1.8e-07 W=4.4e-07 $X=53855 $Y=-39125 $D=0
M89 GND RST 423 GND NM L=1.8e-07 W=4.4e-07 $X=54575 $Y=-42825 $D=0
M90 GND RST 424 GND NM L=1.8e-07 W=4.4e-07 $X=54575 $Y=-39125 $D=0
M91 GND D3 107 GND NM L=1.8e-07 W=2.2e-07 $X=56125 $Y=-26240 $D=0
M92 437 B3 425 GND NM L=1.8e-07 W=4.4e-07 $X=56165 $Y=-17660 $D=0
M93 GND 12 434 GND NM L=1.8e-07 W=2.2e-07 $X=56555 $Y=-42725 $D=0
M94 GND 11 435 GND NM L=1.8e-07 W=2.2e-07 $X=56555 $Y=-39005 $D=0
M95 110 107 GND GND NM L=1.8e-07 W=2.2e-07 $X=56925 $Y=-26240 $D=0
M96 785 462 GND GND NM L=1.8e-07 W=4.4e-07 $X=58535 $Y=-42825 $D=0
M97 786 463 GND GND NM L=1.8e-07 W=4.4e-07 $X=58535 $Y=-39125 $D=0
M98 Q5 CLKREG 785 GND NM L=1.8e-07 W=4.4e-07 $X=58965 $Y=-42825 $D=0
M99 Q4 CLKREG 786 GND NM L=1.8e-07 W=4.4e-07 $X=58965 $Y=-39125 $D=0
M100 GND D4 111 GND NM L=1.8e-07 W=2.2e-07 $X=60585 $Y=-26240 $D=0
M101 464 B4 452 GND NM L=1.8e-07 W=4.4e-07 $X=60625 $Y=-17660 $D=0
M102 787 CLKREG 462 GND NM L=1.8e-07 W=4.4e-07 $X=60905 $Y=-42825 $D=0
M103 788 CLKREG 463 GND NM L=1.8e-07 W=4.4e-07 $X=60905 $Y=-39125 $D=0
M104 GND 476 787 GND NM L=1.8e-07 W=4.4e-07 $X=61335 $Y=-42825 $D=0
M105 GND 477 788 GND NM L=1.8e-07 W=4.4e-07 $X=61335 $Y=-39125 $D=0
M106 114 111 GND GND NM L=1.8e-07 W=2.2e-07 $X=61385 $Y=-26240 $D=0
M107 476 479 GND GND NM L=1.8e-07 W=4.4e-07 $X=62055 $Y=-42825 $D=0
M108 477 480 GND GND NM L=1.8e-07 W=4.4e-07 $X=62055 $Y=-39125 $D=0
M109 GND RST 476 GND NM L=1.8e-07 W=4.4e-07 $X=62775 $Y=-42825 $D=0
M110 GND RST 477 GND NM L=1.8e-07 W=4.4e-07 $X=62775 $Y=-39125 $D=0
M111 GND 14 479 GND NM L=1.8e-07 W=2.2e-07 $X=64755 $Y=-42725 $D=0
M112 GND 13 480 GND NM L=1.8e-07 W=2.2e-07 $X=64755 $Y=-39005 $D=0
M113 GND D5 115 GND NM L=1.8e-07 W=2.2e-07 $X=65045 $Y=-26240 $D=0
M114 491 B5 481 GND NM L=1.8e-07 W=4.4e-07 $X=65085 $Y=-17660 $D=0
M115 118 115 GND GND NM L=1.8e-07 W=2.2e-07 $X=65845 $Y=-26240 $D=0
M116 789 506 GND GND NM L=1.8e-07 W=4.4e-07 $X=66735 $Y=-42825 $D=0
M117 790 507 GND GND NM L=1.8e-07 W=4.4e-07 $X=66735 $Y=-39125 $D=0
M118 Q7 CLKREG 789 GND NM L=1.8e-07 W=4.4e-07 $X=67165 $Y=-42825 $D=0
M119 Q6 CLKREG 790 GND NM L=1.8e-07 W=4.4e-07 $X=67165 $Y=-39125 $D=0
M120 791 CLKREG 506 GND NM L=1.8e-07 W=4.4e-07 $X=69105 $Y=-42825 $D=0
M121 792 CLKREG 507 GND NM L=1.8e-07 W=4.4e-07 $X=69105 $Y=-39125 $D=0
M122 GND D6 119 GND NM L=1.8e-07 W=2.2e-07 $X=69505 $Y=-26240 $D=0
M123 GND 530 791 GND NM L=1.8e-07 W=4.4e-07 $X=69535 $Y=-42825 $D=0
M124 GND 531 792 GND NM L=1.8e-07 W=4.4e-07 $X=69535 $Y=-39125 $D=0
M125 518 B6 508 GND NM L=1.8e-07 W=4.4e-07 $X=69545 $Y=-17660 $D=0
M126 530 532 GND GND NM L=1.8e-07 W=4.4e-07 $X=70255 $Y=-42825 $D=0
M127 531 533 GND GND NM L=1.8e-07 W=4.4e-07 $X=70255 $Y=-39125 $D=0
M128 122 119 GND GND NM L=1.8e-07 W=2.2e-07 $X=70305 $Y=-26240 $D=0
M129 GND RST 530 GND NM L=1.8e-07 W=4.4e-07 $X=70975 $Y=-42825 $D=0
M130 GND RST 531 GND NM L=1.8e-07 W=4.4e-07 $X=70975 $Y=-39125 $D=0
M131 GND 16 532 GND NM L=1.8e-07 W=2.2e-07 $X=72955 $Y=-42725 $D=0
M132 GND 15 533 GND NM L=1.8e-07 W=2.2e-07 $X=72955 $Y=-39005 $D=0
M133 GND D7 124 GND NM L=1.8e-07 W=2.2e-07 $X=73965 $Y=-26240 $D=0
M134 545 B7 535 GND NM L=1.8e-07 W=4.4e-07 $X=74005 $Y=-17660 $D=0
M135 127 124 GND GND NM L=1.8e-07 W=2.2e-07 $X=74765 $Y=-26240 $D=0
M136 793 559 GND GND NM L=1.8e-07 W=4.4e-07 $X=74935 $Y=-42825 $D=0
M137 794 560 GND GND NM L=1.8e-07 W=4.4e-07 $X=74935 $Y=-39125 $D=0
M138 Q9 CLKREG 793 GND NM L=1.8e-07 W=4.4e-07 $X=75365 $Y=-42825 $D=0
M139 Q8 CLKREG 794 GND NM L=1.8e-07 W=4.4e-07 $X=75365 $Y=-39125 $D=0
M140 795 CLKREG 559 GND NM L=1.8e-07 W=4.4e-07 $X=77305 $Y=-42825 $D=0
M141 796 CLKREG 560 GND NM L=1.8e-07 W=4.4e-07 $X=77305 $Y=-39125 $D=0
M142 GND 582 795 GND NM L=1.8e-07 W=4.4e-07 $X=77735 $Y=-42825 $D=0
M143 GND 583 796 GND NM L=1.8e-07 W=4.4e-07 $X=77735 $Y=-39125 $D=0
M144 GND D8 128 GND NM L=1.8e-07 W=2.2e-07 $X=78425 $Y=-26240 $D=0
M145 582 586 GND GND NM L=1.8e-07 W=4.4e-07 $X=78455 $Y=-42825 $D=0
M146 583 587 GND GND NM L=1.8e-07 W=4.4e-07 $X=78455 $Y=-39125 $D=0
M147 572 B8 562 GND NM L=1.8e-07 W=4.4e-07 $X=78465 $Y=-17660 $D=0
M148 GND RST 582 GND NM L=1.8e-07 W=4.4e-07 $X=79175 $Y=-42825 $D=0
M149 GND RST 583 GND NM L=1.8e-07 W=4.4e-07 $X=79175 $Y=-39125 $D=0
M150 131 128 GND GND NM L=1.8e-07 W=2.2e-07 $X=79225 $Y=-26240 $D=0
M151 GND 18 586 GND NM L=1.8e-07 W=2.2e-07 $X=81155 $Y=-42725 $D=0
M152 GND 17 587 GND NM L=1.8e-07 W=2.2e-07 $X=81155 $Y=-39005 $D=0
M153 GND D9 132 GND NM L=1.8e-07 W=2.2e-07 $X=82885 $Y=-26240 $D=0
M154 599 B9 589 GND NM L=1.8e-07 W=4.4e-07 $X=82925 $Y=-17660 $D=0
M155 797 613 GND GND NM L=1.8e-07 W=4.4e-07 $X=83135 $Y=-42825 $D=0
M156 798 614 GND GND NM L=1.8e-07 W=4.4e-07 $X=83135 $Y=-39125 $D=0
M157 Q11 CLKREG 797 GND NM L=1.8e-07 W=4.4e-07 $X=83565 $Y=-42825 $D=0
M158 Q10 CLKREG 798 GND NM L=1.8e-07 W=4.4e-07 $X=83565 $Y=-39125 $D=0
M159 135 132 GND GND NM L=1.8e-07 W=2.2e-07 $X=83685 $Y=-26240 $D=0
M160 799 CLKREG 613 GND NM L=1.8e-07 W=4.4e-07 $X=85505 $Y=-42825 $D=0
M161 800 CLKREG 614 GND NM L=1.8e-07 W=4.4e-07 $X=85505 $Y=-39125 $D=0
M162 GND 627 799 GND NM L=1.8e-07 W=4.4e-07 $X=85935 $Y=-42825 $D=0
M163 GND 628 800 GND NM L=1.8e-07 W=4.4e-07 $X=85935 $Y=-39125 $D=0
M164 627 639 GND GND NM L=1.8e-07 W=4.4e-07 $X=86655 $Y=-42825 $D=0
M165 628 640 GND GND NM L=1.8e-07 W=4.4e-07 $X=86655 $Y=-39125 $D=0
M166 GND D10 136 GND NM L=1.8e-07 W=2.2e-07 $X=87345 $Y=-26240 $D=0
M167 GND RST 627 GND NM L=1.8e-07 W=4.4e-07 $X=87375 $Y=-42825 $D=0
M168 GND RST 628 GND NM L=1.8e-07 W=4.4e-07 $X=87375 $Y=-39125 $D=0
M169 626 B10 616 GND NM L=1.8e-07 W=4.4e-07 $X=87385 $Y=-17660 $D=0
M170 139 136 GND GND NM L=1.8e-07 W=2.2e-07 $X=88145 $Y=-26240 $D=0
M171 GND 20 639 GND NM L=1.8e-07 W=2.2e-07 $X=89355 $Y=-42725 $D=0
M172 GND 19 640 GND NM L=1.8e-07 W=2.2e-07 $X=89355 $Y=-39005 $D=0
M173 801 667 GND GND NM L=1.8e-07 W=4.4e-07 $X=91335 $Y=-42825 $D=0
M174 802 668 GND GND NM L=1.8e-07 W=4.4e-07 $X=91335 $Y=-39125 $D=0
M175 Q13 CLKREG 801 GND NM L=1.8e-07 W=4.4e-07 $X=91765 $Y=-42825 $D=0
M176 Q12 CLKREG 802 GND NM L=1.8e-07 W=4.4e-07 $X=91765 $Y=-39125 $D=0
M177 GND D11 140 GND NM L=1.8e-07 W=2.2e-07 $X=91805 $Y=-26240 $D=0
M178 655 B11 643 GND NM L=1.8e-07 W=4.4e-07 $X=91845 $Y=-17660 $D=0
M179 143 140 GND GND NM L=1.8e-07 W=2.2e-07 $X=92605 $Y=-26240 $D=0
M180 803 CLKREG 667 GND NM L=1.8e-07 W=4.4e-07 $X=93705 $Y=-42825 $D=0
M181 804 CLKREG 668 GND NM L=1.8e-07 W=4.4e-07 $X=93705 $Y=-39125 $D=0
M182 GND 671 803 GND NM L=1.8e-07 W=4.4e-07 $X=94135 $Y=-42825 $D=0
M183 GND 672 804 GND NM L=1.8e-07 W=4.4e-07 $X=94135 $Y=-39125 $D=0
M184 671 683 GND GND NM L=1.8e-07 W=4.4e-07 $X=94855 $Y=-42825 $D=0
M185 672 684 GND GND NM L=1.8e-07 W=4.4e-07 $X=94855 $Y=-39125 $D=0
M186 GND RST 671 GND NM L=1.8e-07 W=4.4e-07 $X=95575 $Y=-42825 $D=0
M187 GND RST 672 GND NM L=1.8e-07 W=4.4e-07 $X=95575 $Y=-39125 $D=0
M188 GND D12 144 GND NM L=1.8e-07 W=2.2e-07 $X=96265 $Y=-26240 $D=0
M189 682 B12 670 GND NM L=1.8e-07 W=4.4e-07 $X=96305 $Y=-17660 $D=0
M190 147 144 GND GND NM L=1.8e-07 W=2.2e-07 $X=97065 $Y=-26240 $D=0
M191 GND 22 683 GND NM L=1.8e-07 W=2.2e-07 $X=97555 $Y=-42725 $D=0
M192 GND 21 684 GND NM L=1.8e-07 W=2.2e-07 $X=97555 $Y=-39005 $D=0
M193 805 719 GND GND NM L=1.8e-07 W=4.4e-07 $X=99535 $Y=-42825 $D=0
M194 806 720 GND GND NM L=1.8e-07 W=4.4e-07 $X=99535 $Y=-39125 $D=0
M195 Q15 CLKREG 805 GND NM L=1.8e-07 W=4.4e-07 $X=99965 $Y=-42825 $D=0
M196 Q14 CLKREG 806 GND NM L=1.8e-07 W=4.4e-07 $X=99965 $Y=-39125 $D=0
M197 GND D13 148 GND NM L=1.8e-07 W=2.2e-07 $X=100725 $Y=-26240 $D=0
M198 709 B13 699 GND NM L=1.8e-07 W=4.4e-07 $X=100765 $Y=-17660 $D=0
M199 151 148 GND GND NM L=1.8e-07 W=2.2e-07 $X=101525 $Y=-26240 $D=0
M200 807 CLKREG 719 GND NM L=1.8e-07 W=4.4e-07 $X=101905 $Y=-42825 $D=0
M201 808 CLKREG 720 GND NM L=1.8e-07 W=4.4e-07 $X=101905 $Y=-39125 $D=0
M202 GND 724 807 GND NM L=1.8e-07 W=4.4e-07 $X=102335 $Y=-42825 $D=0
M203 GND 725 808 GND NM L=1.8e-07 W=4.4e-07 $X=102335 $Y=-39125 $D=0
M204 724 736 GND GND NM L=1.8e-07 W=4.4e-07 $X=103055 $Y=-42825 $D=0
M205 725 737 GND GND NM L=1.8e-07 W=4.4e-07 $X=103055 $Y=-39125 $D=0
M206 GND RST 724 GND NM L=1.8e-07 W=4.4e-07 $X=103775 $Y=-42825 $D=0
M207 GND RST 725 GND NM L=1.8e-07 W=4.4e-07 $X=103775 $Y=-39125 $D=0
M208 GND D14 152 GND NM L=1.8e-07 W=2.2e-07 $X=105185 $Y=-26240 $D=0
M209 738 B14 726 GND NM L=1.8e-07 W=4.4e-07 $X=105225 $Y=-17660 $D=0
M210 GND 24 736 GND NM L=1.8e-07 W=2.2e-07 $X=105755 $Y=-42725 $D=0
M211 GND 23 737 GND NM L=1.8e-07 W=2.2e-07 $X=105755 $Y=-39005 $D=0
M212 155 152 GND GND NM L=1.8e-07 W=2.2e-07 $X=105985 $Y=-26240 $D=0
M213 GND D15 156 GND NM L=1.8e-07 W=2.2e-07 $X=109645 $Y=-26240 $D=0
M214 761 B15 751 GND NM L=1.8e-07 W=4.4e-07 $X=109685 $Y=-17660 $D=0
M215 159 156 GND GND NM L=1.8e-07 W=2.2e-07 $X=110445 $Y=-26240 $D=0
M216 823 28 31 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=-840 $D=4
M217 VDD 29 824 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=20 $D=4
M218 825 28 34 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=2780 $D=4
M219 826 30 825 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=3210 $D=4
M220 VDD A0 826 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=3640 $D=4
M221 827 28 35 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=6400 $D=4
M222 828 A1 827 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=6830 $D=4
M223 VDD 29 828 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=7260 $D=4
M224 VDD A0 829 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=10880 $D=4
M225 831 A1 830 VDD PM L=1.8e-07 W=1.32e-06 $X=-9375 $Y=21310 $D=4
M226 194 31 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=-7840 $D=4
M227 195 34 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=-3200 $D=4
M228 196 35 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=1440 $D=4
M229 197 36 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=6080 $D=4
M230 198 37 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=10720 $D=4
M231 VDD 199 4 VDD PM L=1.8e-07 W=4.4e-07 $X=-6575 $Y=13420 $D=4
M232 199 38 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=15360 $D=4
M233 VDD 200 3 VDD PM L=1.8e-07 W=4.4e-07 $X=-6575 $Y=18060 $D=4
M234 200 32 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=20000 $D=4
M235 VDD CLK 200 VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=20720 $D=4
M236 201 33 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=24640 $D=4
M237 VDD CLK 201 VDD PM L=1.8e-07 W=8.8e-07 $X=-6575 $Y=25360 $D=4
M238 VDD 42 287 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=-13910 $D=4
M239 VDD 43 288 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=-11550 $D=4
M240 VDD 44 289 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=1330 $D=4
M241 VDD 45 290 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=3690 $D=4
M242 VDD 46 291 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=16570 $D=4
M243 VDD 47 292 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=18930 $D=4
M244 VDD 48 293 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=31810 $D=4
M245 VDD 49 294 VDD PM L=1.8e-07 W=8.8e-07 $X=20415 $Y=34170 $D=4
M246 VDD 296 306 VDD PM L=1.8e-07 W=8.8e-07 $X=23195 $Y=47050 $D=4
M247 VDD 298 308 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=-13910 $D=4
M248 VDD 299 309 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=-11550 $D=4
M249 VDD 300 310 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=1330 $D=4
M250 VDD 301 311 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=3690 $D=4
M251 VDD 302 312 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=16570 $D=4
M252 VDD 303 313 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=18930 $D=4
M253 VDD 304 314 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=31810 $D=4
M254 VDD 305 315 VDD PM L=1.8e-07 W=8.8e-07 $X=25055 $Y=34170 $D=4
M255 307 297 VDD VDD PM L=1.8e-07 W=1.76e-06 $X=25935 $Y=-30030 $D=4
M256 54 GND VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27155 $Y=-26790 $D=4
M257 325 324 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29855 $Y=-28710 $D=4
M258 40 52 832 VDD PM L=1.8e-07 W=8.8e-07 $X=31585 $Y=-26790 $D=4
M259 833 54 40 VDD PM L=1.8e-07 W=8.8e-07 $X=32305 $Y=-26790 $D=4
M260 834 55 41 VDD PM L=1.8e-07 W=8.8e-07 $X=32305 $Y=47050 $D=4
M261 VDD 325 326 VDD PM L=1.8e-07 W=8.8e-07 $X=32555 $Y=-29150 $D=4
M262 VDD 64 833 VDD PM L=1.8e-07 W=8.8e-07 $X=32735 $Y=-26790 $D=4
M263 VDD 65 834 VDD PM L=1.8e-07 W=8.8e-07 $X=32735 $Y=47050 $D=4
M264 835 66 ADD7 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=-13910 $D=4
M265 836 67 ADD6 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=-11550 $D=4
M266 837 68 ADD5 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=1330 $D=4
M267 838 69 ADD4 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=3690 $D=4
M268 839 70 ADD3 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=16570 $D=4
M269 840 71 ADD2 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=18930 $D=4
M270 841 72 ADD1 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=31810 $D=4
M271 842 73 ADD0 VDD PM L=1.8e-07 W=8.8e-07 $X=36185 $Y=34170 $D=4
M272 VDD 77 835 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=-13910 $D=4
M273 VDD 78 836 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=-11550 $D=4
M274 VDD 79 837 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=1330 $D=4
M275 VDD 80 838 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=3690 $D=4
M276 VDD 81 839 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=16570 $D=4
M277 VDD 82 840 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=18930 $D=4
M278 VDD 83 841 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=31810 $D=4
M279 VDD 84 842 VDD PM L=1.8e-07 W=8.8e-07 $X=36615 $Y=34170 $D=4
M280 Q1 365 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42135 $Y=-46270 $D=4
M281 Q0 366 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42135 $Y=-36120 $D=4
M282 VDD D0 94 VDD PM L=1.8e-07 W=4.4e-07 $X=42785 $Y=-24530 $D=4
M283 VDD 342 342 VDD PM L=1.8e-07 W=3.3e-06 $X=42785 $Y=-15250 $D=4
M284 98 94 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=43505 $Y=-24530 $D=4
M285 VDD CLKREG 365 VDD PM L=1.8e-07 W=8.8e-07 $X=44835 $Y=-46270 $D=4
M286 VDD CLKREG 366 VDD PM L=1.8e-07 W=8.8e-07 $X=44835 $Y=-36120 $D=4
M287 843 382 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=45555 $Y=-46270 $D=4
M288 844 383 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=45555 $Y=-36120 $D=4
M289 845 RST 843 VDD PM L=1.8e-07 W=8.8e-07 $X=45985 $Y=-46270 $D=4
M290 846 RST 844 VDD PM L=1.8e-07 W=8.8e-07 $X=45985 $Y=-36120 $D=4
M291 369 CLKREG 845 VDD PM L=1.8e-07 W=8.8e-07 $X=46415 $Y=-46270 $D=4
M292 370 CLKREG 846 VDD PM L=1.8e-07 W=8.8e-07 $X=46415 $Y=-36120 $D=4
M293 VDD D1 99 VDD PM L=1.8e-07 W=4.4e-07 $X=47245 $Y=-24530 $D=4
M294 VDD 371 371 VDD PM L=1.8e-07 W=3.3e-06 $X=47245 $Y=-15250 $D=4
M295 102 99 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=47965 $Y=-24530 $D=4
M296 VDD 10 382 VDD PM L=1.8e-07 W=4.4e-07 $X=48355 $Y=-46270 $D=4
M297 VDD 9 383 VDD PM L=1.8e-07 W=4.4e-07 $X=48355 $Y=-35680 $D=4
M298 Q3 409 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50335 $Y=-46270 $D=4
M299 Q2 410 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50335 $Y=-36120 $D=4
M300 VDD D2 103 VDD PM L=1.8e-07 W=4.4e-07 $X=51705 $Y=-24530 $D=4
M301 VDD 398 398 VDD PM L=1.8e-07 W=3.3e-06 $X=51705 $Y=-15250 $D=4
M302 106 103 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=52425 $Y=-24530 $D=4
M303 VDD CLKREG 409 VDD PM L=1.8e-07 W=8.8e-07 $X=53035 $Y=-46270 $D=4
M304 VDD CLKREG 410 VDD PM L=1.8e-07 W=8.8e-07 $X=53035 $Y=-36120 $D=4
M305 847 434 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53755 $Y=-46270 $D=4
M306 848 435 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53755 $Y=-36120 $D=4
M307 849 RST 847 VDD PM L=1.8e-07 W=8.8e-07 $X=54185 $Y=-46270 $D=4
M308 850 RST 848 VDD PM L=1.8e-07 W=8.8e-07 $X=54185 $Y=-36120 $D=4
M309 423 CLKREG 849 VDD PM L=1.8e-07 W=8.8e-07 $X=54615 $Y=-46270 $D=4
M310 424 CLKREG 850 VDD PM L=1.8e-07 W=8.8e-07 $X=54615 $Y=-36120 $D=4
M311 VDD D3 107 VDD PM L=1.8e-07 W=4.4e-07 $X=56165 $Y=-24530 $D=4
M312 VDD 425 425 VDD PM L=1.8e-07 W=3.3e-06 $X=56165 $Y=-15250 $D=4
M313 VDD 12 434 VDD PM L=1.8e-07 W=4.4e-07 $X=56555 $Y=-46270 $D=4
M314 VDD 11 435 VDD PM L=1.8e-07 W=4.4e-07 $X=56555 $Y=-35680 $D=4
M315 110 107 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=56885 $Y=-24530 $D=4
M316 Q5 462 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=58535 $Y=-46270 $D=4
M317 Q4 463 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=58535 $Y=-36120 $D=4
M318 VDD D4 111 VDD PM L=1.8e-07 W=4.4e-07 $X=60625 $Y=-24530 $D=4
M319 VDD 452 452 VDD PM L=1.8e-07 W=3.3e-06 $X=60625 $Y=-15250 $D=4
M320 VDD CLKREG 462 VDD PM L=1.8e-07 W=8.8e-07 $X=61235 $Y=-46270 $D=4
M321 VDD CLKREG 463 VDD PM L=1.8e-07 W=8.8e-07 $X=61235 $Y=-36120 $D=4
M322 114 111 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=61345 $Y=-24530 $D=4
M323 851 479 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61955 $Y=-46270 $D=4
M324 852 480 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61955 $Y=-36120 $D=4
M325 853 RST 851 VDD PM L=1.8e-07 W=8.8e-07 $X=62385 $Y=-46270 $D=4
M326 854 RST 852 VDD PM L=1.8e-07 W=8.8e-07 $X=62385 $Y=-36120 $D=4
M327 476 CLKREG 853 VDD PM L=1.8e-07 W=8.8e-07 $X=62815 $Y=-46270 $D=4
M328 477 CLKREG 854 VDD PM L=1.8e-07 W=8.8e-07 $X=62815 $Y=-36120 $D=4
M329 VDD 14 479 VDD PM L=1.8e-07 W=4.4e-07 $X=64755 $Y=-46270 $D=4
M330 VDD 13 480 VDD PM L=1.8e-07 W=4.4e-07 $X=64755 $Y=-35680 $D=4
M331 VDD D5 115 VDD PM L=1.8e-07 W=4.4e-07 $X=65085 $Y=-24530 $D=4
M332 VDD 481 481 VDD PM L=1.8e-07 W=3.3e-06 $X=65085 $Y=-15250 $D=4
M333 118 115 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=65805 $Y=-24530 $D=4
M334 Q7 506 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=66735 $Y=-46270 $D=4
M335 Q6 507 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=66735 $Y=-36120 $D=4
M336 VDD CLKREG 506 VDD PM L=1.8e-07 W=8.8e-07 $X=69435 $Y=-46270 $D=4
M337 VDD CLKREG 507 VDD PM L=1.8e-07 W=8.8e-07 $X=69435 $Y=-36120 $D=4
M338 VDD D6 119 VDD PM L=1.8e-07 W=4.4e-07 $X=69545 $Y=-24530 $D=4
M339 VDD 508 508 VDD PM L=1.8e-07 W=3.3e-06 $X=69545 $Y=-15250 $D=4
M340 855 532 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=70155 $Y=-46270 $D=4
M341 856 533 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=70155 $Y=-36120 $D=4
M342 122 119 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=70265 $Y=-24530 $D=4
M343 857 RST 855 VDD PM L=1.8e-07 W=8.8e-07 $X=70585 $Y=-46270 $D=4
M344 858 RST 856 VDD PM L=1.8e-07 W=8.8e-07 $X=70585 $Y=-36120 $D=4
M345 530 CLKREG 857 VDD PM L=1.8e-07 W=8.8e-07 $X=71015 $Y=-46270 $D=4
M346 531 CLKREG 858 VDD PM L=1.8e-07 W=8.8e-07 $X=71015 $Y=-36120 $D=4
M347 VDD 16 532 VDD PM L=1.8e-07 W=4.4e-07 $X=72955 $Y=-46270 $D=4
M348 VDD 15 533 VDD PM L=1.8e-07 W=4.4e-07 $X=72955 $Y=-35680 $D=4
M349 VDD D7 124 VDD PM L=1.8e-07 W=4.4e-07 $X=74005 $Y=-24530 $D=4
M350 VDD 535 535 VDD PM L=1.8e-07 W=3.3e-06 $X=74005 $Y=-15250 $D=4
M351 127 124 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=74725 $Y=-24530 $D=4
M352 Q9 559 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=74935 $Y=-46270 $D=4
M353 Q8 560 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=74935 $Y=-36120 $D=4
M354 VDD CLKREG 559 VDD PM L=1.8e-07 W=8.8e-07 $X=77635 $Y=-46270 $D=4
M355 VDD CLKREG 560 VDD PM L=1.8e-07 W=8.8e-07 $X=77635 $Y=-36120 $D=4
M356 859 586 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=78355 $Y=-46270 $D=4
M357 860 587 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=78355 $Y=-36120 $D=4
M358 VDD D8 128 VDD PM L=1.8e-07 W=4.4e-07 $X=78465 $Y=-24530 $D=4
M359 VDD 562 562 VDD PM L=1.8e-07 W=3.3e-06 $X=78465 $Y=-15250 $D=4
M360 861 RST 859 VDD PM L=1.8e-07 W=8.8e-07 $X=78785 $Y=-46270 $D=4
M361 862 RST 860 VDD PM L=1.8e-07 W=8.8e-07 $X=78785 $Y=-36120 $D=4
M362 131 128 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=79185 $Y=-24530 $D=4
M363 582 CLKREG 861 VDD PM L=1.8e-07 W=8.8e-07 $X=79215 $Y=-46270 $D=4
M364 583 CLKREG 862 VDD PM L=1.8e-07 W=8.8e-07 $X=79215 $Y=-36120 $D=4
M365 VDD 18 586 VDD PM L=1.8e-07 W=4.4e-07 $X=81155 $Y=-46270 $D=4
M366 VDD 17 587 VDD PM L=1.8e-07 W=4.4e-07 $X=81155 $Y=-35680 $D=4
M367 VDD D9 132 VDD PM L=1.8e-07 W=4.4e-07 $X=82925 $Y=-24530 $D=4
M368 VDD 589 589 VDD PM L=1.8e-07 W=3.3e-06 $X=82925 $Y=-15250 $D=4
M369 Q11 613 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=83135 $Y=-46270 $D=4
M370 Q10 614 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=83135 $Y=-36120 $D=4
M371 135 132 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=83645 $Y=-24530 $D=4
M372 VDD CLKREG 613 VDD PM L=1.8e-07 W=8.8e-07 $X=85835 $Y=-46270 $D=4
M373 VDD CLKREG 614 VDD PM L=1.8e-07 W=8.8e-07 $X=85835 $Y=-36120 $D=4
M374 863 639 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=86555 $Y=-46270 $D=4
M375 864 640 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=86555 $Y=-36120 $D=4
M376 865 RST 863 VDD PM L=1.8e-07 W=8.8e-07 $X=86985 $Y=-46270 $D=4
M377 866 RST 864 VDD PM L=1.8e-07 W=8.8e-07 $X=86985 $Y=-36120 $D=4
M378 VDD D10 136 VDD PM L=1.8e-07 W=4.4e-07 $X=87385 $Y=-24530 $D=4
M379 VDD 616 616 VDD PM L=1.8e-07 W=3.3e-06 $X=87385 $Y=-15250 $D=4
M380 627 CLKREG 865 VDD PM L=1.8e-07 W=8.8e-07 $X=87415 $Y=-46270 $D=4
M381 628 CLKREG 866 VDD PM L=1.8e-07 W=8.8e-07 $X=87415 $Y=-36120 $D=4
M382 139 136 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=88105 $Y=-24530 $D=4
M383 VDD 20 639 VDD PM L=1.8e-07 W=4.4e-07 $X=89355 $Y=-46270 $D=4
M384 VDD 19 640 VDD PM L=1.8e-07 W=4.4e-07 $X=89355 $Y=-35680 $D=4
M385 Q13 667 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=91335 $Y=-46270 $D=4
M386 Q12 668 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=91335 $Y=-36120 $D=4
M387 VDD D11 140 VDD PM L=1.8e-07 W=4.4e-07 $X=91845 $Y=-24530 $D=4
M388 VDD 643 643 VDD PM L=1.8e-07 W=3.3e-06 $X=91845 $Y=-15250 $D=4
M389 143 140 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=92565 $Y=-24530 $D=4
M390 VDD CLKREG 667 VDD PM L=1.8e-07 W=8.8e-07 $X=94035 $Y=-46270 $D=4
M391 VDD CLKREG 668 VDD PM L=1.8e-07 W=8.8e-07 $X=94035 $Y=-36120 $D=4
M392 867 683 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=94755 $Y=-46270 $D=4
M393 868 684 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=94755 $Y=-36120 $D=4
M394 869 RST 867 VDD PM L=1.8e-07 W=8.8e-07 $X=95185 $Y=-46270 $D=4
M395 870 RST 868 VDD PM L=1.8e-07 W=8.8e-07 $X=95185 $Y=-36120 $D=4
M396 671 CLKREG 869 VDD PM L=1.8e-07 W=8.8e-07 $X=95615 $Y=-46270 $D=4
M397 672 CLKREG 870 VDD PM L=1.8e-07 W=8.8e-07 $X=95615 $Y=-36120 $D=4
M398 VDD D12 144 VDD PM L=1.8e-07 W=4.4e-07 $X=96305 $Y=-24530 $D=4
M399 VDD 670 670 VDD PM L=1.8e-07 W=3.3e-06 $X=96305 $Y=-15250 $D=4
M400 147 144 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=97025 $Y=-24530 $D=4
M401 VDD 22 683 VDD PM L=1.8e-07 W=4.4e-07 $X=97555 $Y=-46270 $D=4
M402 VDD 21 684 VDD PM L=1.8e-07 W=4.4e-07 $X=97555 $Y=-35680 $D=4
M403 Q15 719 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=99535 $Y=-46270 $D=4
M404 Q14 720 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=99535 $Y=-36120 $D=4
M405 VDD D13 148 VDD PM L=1.8e-07 W=4.4e-07 $X=100765 $Y=-24530 $D=4
M406 VDD 699 699 VDD PM L=1.8e-07 W=3.3e-06 $X=100765 $Y=-15250 $D=4
M407 151 148 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=101485 $Y=-24530 $D=4
M408 VDD CLKREG 719 VDD PM L=1.8e-07 W=8.8e-07 $X=102235 $Y=-46270 $D=4
M409 VDD CLKREG 720 VDD PM L=1.8e-07 W=8.8e-07 $X=102235 $Y=-36120 $D=4
M410 871 736 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=102955 $Y=-46270 $D=4
M411 872 737 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=102955 $Y=-36120 $D=4
M412 873 RST 871 VDD PM L=1.8e-07 W=8.8e-07 $X=103385 $Y=-46270 $D=4
M413 874 RST 872 VDD PM L=1.8e-07 W=8.8e-07 $X=103385 $Y=-36120 $D=4
M414 724 CLKREG 873 VDD PM L=1.8e-07 W=8.8e-07 $X=103815 $Y=-46270 $D=4
M415 725 CLKREG 874 VDD PM L=1.8e-07 W=8.8e-07 $X=103815 $Y=-36120 $D=4
M416 VDD D14 152 VDD PM L=1.8e-07 W=4.4e-07 $X=105225 $Y=-24530 $D=4
M417 VDD 726 726 VDD PM L=1.8e-07 W=3.3e-06 $X=105225 $Y=-15250 $D=4
M418 VDD 24 736 VDD PM L=1.8e-07 W=4.4e-07 $X=105755 $Y=-46270 $D=4
M419 VDD 23 737 VDD PM L=1.8e-07 W=4.4e-07 $X=105755 $Y=-35680 $D=4
M420 155 152 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=105945 $Y=-24530 $D=4
M421 VDD D15 156 VDD PM L=1.8e-07 W=4.4e-07 $X=109685 $Y=-24530 $D=4
M422 VDD 751 751 VDD PM L=1.8e-07 W=3.3e-06 $X=109685 $Y=-15250 $D=4
M423 159 156 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=110405 $Y=-24530 $D=4
X424 GND 364 354 INVB0 n18_CDNS_6738713766025 $T=43685 -17660 1 180 $X=42845 $Y=-18010
X425 GND 393 381 INVB1 n18_CDNS_6738713766025 $T=48145 -17660 1 180 $X=47305 $Y=-18010
X426 GND 420 408 INVB2 n18_CDNS_6738713766025 $T=52605 -17660 1 180 $X=51765 $Y=-18010
X427 GND 447 437 INVB3 n18_CDNS_6738713766025 $T=57065 -17660 1 180 $X=56225 $Y=-18010
X428 GND 474 464 INVB4 n18_CDNS_6738713766025 $T=61525 -17660 1 180 $X=60685 $Y=-18010
X429 GND 501 491 INVB5 n18_CDNS_6738713766025 $T=65985 -17660 1 180 $X=65145 $Y=-18010
X430 GND 528 518 INVB6 n18_CDNS_6738713766025 $T=70445 -17660 1 180 $X=69605 $Y=-18010
X431 GND 555 545 INVB7 n18_CDNS_6738713766025 $T=74905 -17660 1 180 $X=74065 $Y=-18010
X432 GND 584 572 INVB8 n18_CDNS_6738713766025 $T=79365 -17660 1 180 $X=78525 $Y=-18010
X433 GND 611 599 INVB9 n18_CDNS_6738713766025 $T=83825 -17660 1 180 $X=82985 $Y=-18010
X434 GND 638 626 INVB10 n18_CDNS_6738713766025 $T=88285 -17660 1 180 $X=87445 $Y=-18010
X435 GND 665 655 INVB11 n18_CDNS_6738713766025 $T=92745 -17660 1 180 $X=91905 $Y=-18010
X436 GND 694 682 INVB12 n18_CDNS_6738713766025 $T=97205 -17660 1 180 $X=96365 $Y=-18010
X437 GND 721 709 INVB13 n18_CDNS_6738713766025 $T=101665 -17660 1 180 $X=100825 $Y=-18010
X438 GND 748 738 INVB14 n18_CDNS_6738713766025 $T=106125 -17660 1 180 $X=105285 $Y=-18010
X439 GND 771 761 INVB15 n18_CDNS_6738713766025 $T=110585 -17660 1 180 $X=109745 $Y=-18010
X440 VDD 364 342 p18_CDNS_6738713766022 $T=43685 -15250 1 180 $X=42595 $Y=-15680
X441 VDD 393 371 p18_CDNS_6738713766022 $T=48145 -15250 1 180 $X=47055 $Y=-15680
X442 VDD 420 398 p18_CDNS_6738713766022 $T=52605 -15250 1 180 $X=51515 $Y=-15680
X443 VDD 447 425 p18_CDNS_6738713766022 $T=57065 -15250 1 180 $X=55975 $Y=-15680
X444 VDD 474 452 p18_CDNS_6738713766022 $T=61525 -15250 1 180 $X=60435 $Y=-15680
X445 VDD 501 481 p18_CDNS_6738713766022 $T=65985 -15250 1 180 $X=64895 $Y=-15680
X446 VDD 528 508 p18_CDNS_6738713766022 $T=70445 -15250 1 180 $X=69355 $Y=-15680
X447 VDD 555 535 p18_CDNS_6738713766022 $T=74905 -15250 1 180 $X=73815 $Y=-15680
X448 VDD 584 562 p18_CDNS_6738713766022 $T=79365 -15250 1 180 $X=78275 $Y=-15680
X449 VDD 611 589 p18_CDNS_6738713766022 $T=83825 -15250 1 180 $X=82735 $Y=-15680
X450 VDD 638 616 p18_CDNS_6738713766022 $T=88285 -15250 1 180 $X=87195 $Y=-15680
X451 VDD 665 643 p18_CDNS_6738713766022 $T=92745 -15250 1 180 $X=91655 $Y=-15680
X452 VDD 694 670 p18_CDNS_6738713766022 $T=97205 -15250 1 180 $X=96115 $Y=-15680
X453 VDD 721 699 p18_CDNS_6738713766022 $T=101665 -15250 1 180 $X=100575 $Y=-15680
X454 VDD 748 726 p18_CDNS_6738713766022 $T=106125 -15250 1 180 $X=105035 $Y=-15680
X455 VDD 771 751 p18_CDNS_6738713766022 $T=110585 -15250 1 180 $X=109495 $Y=-15680
X456 B0 INVB0 PCEN VDD p18_CDNS_6738713766029 $T=43015 38420 0 270 $X=42585 $Y=37330
X457 B1 INVB1 PCEN VDD p18_CDNS_6738713766029 $T=47475 38420 0 270 $X=47045 $Y=37330
X458 B2 INVB2 PCEN VDD p18_CDNS_6738713766029 $T=51935 38420 0 270 $X=51505 $Y=37330
X459 B3 INVB3 PCEN VDD p18_CDNS_6738713766029 $T=56395 38420 0 270 $X=55965 $Y=37330
X460 B4 INVB4 PCEN VDD p18_CDNS_6738713766029 $T=60855 38420 0 270 $X=60425 $Y=37330
X461 B5 INVB5 PCEN VDD p18_CDNS_6738713766029 $T=65315 38420 0 270 $X=64885 $Y=37330
X462 B6 INVB6 PCEN VDD p18_CDNS_6738713766029 $T=69775 38420 0 270 $X=69345 $Y=37330
X463 B7 INVB7 PCEN VDD p18_CDNS_6738713766029 $T=74235 38420 0 270 $X=73805 $Y=37330
X464 B8 INVB8 PCEN VDD p18_CDNS_6738713766029 $T=78695 38420 0 270 $X=78265 $Y=37330
X465 B9 INVB9 PCEN VDD p18_CDNS_6738713766029 $T=83155 38420 0 270 $X=82725 $Y=37330
X466 B10 INVB10 PCEN VDD p18_CDNS_6738713766029 $T=87615 38420 0 270 $X=87185 $Y=37330
X467 B11 INVB11 PCEN VDD p18_CDNS_6738713766029 $T=92075 38420 0 270 $X=91645 $Y=37330
X468 B12 INVB12 PCEN VDD p18_CDNS_6738713766029 $T=96535 38420 0 270 $X=96105 $Y=37330
X469 B13 INVB13 PCEN VDD p18_CDNS_6738713766029 $T=100995 38420 0 270 $X=100565 $Y=37330
X470 B14 INVB14 PCEN VDD p18_CDNS_6738713766029 $T=105455 38420 0 270 $X=105025 $Y=37330
X471 B15 INVB15 PCEN VDD p18_CDNS_6738713766029 $T=109915 38420 0 270 $X=109485 $Y=37330
X472 GND 354 SAEN n18_CDNS_6738713766021 $T=42795 -19290 1 90 $X=42445 $Y=-19950
X473 GND 381 SAEN n18_CDNS_6738713766021 $T=47255 -19290 1 90 $X=46905 $Y=-19950
X474 GND 408 SAEN n18_CDNS_6738713766021 $T=51715 -19290 1 90 $X=51365 $Y=-19950
X475 GND 437 SAEN n18_CDNS_6738713766021 $T=56175 -19290 1 90 $X=55825 $Y=-19950
X476 GND 464 SAEN n18_CDNS_6738713766021 $T=60635 -19290 1 90 $X=60285 $Y=-19950
X477 GND 491 SAEN n18_CDNS_6738713766021 $T=65095 -19290 1 90 $X=64745 $Y=-19950
X478 GND 518 SAEN n18_CDNS_6738713766021 $T=69555 -19290 1 90 $X=69205 $Y=-19950
X479 GND 545 SAEN n18_CDNS_6738713766021 $T=74015 -19290 1 90 $X=73665 $Y=-19950
X480 GND 572 SAEN n18_CDNS_6738713766021 $T=78475 -19290 1 90 $X=78125 $Y=-19950
X481 GND 599 SAEN n18_CDNS_6738713766021 $T=82935 -19290 1 90 $X=82585 $Y=-19950
X482 GND 626 SAEN n18_CDNS_6738713766021 $T=87395 -19290 1 90 $X=87045 $Y=-19950
X483 GND 655 SAEN n18_CDNS_6738713766021 $T=91855 -19290 1 90 $X=91505 $Y=-19950
X484 GND 682 SAEN n18_CDNS_6738713766021 $T=96315 -19290 1 90 $X=95965 $Y=-19950
X485 GND 709 SAEN n18_CDNS_6738713766021 $T=100775 -19290 1 90 $X=100425 $Y=-19950
X486 GND 738 SAEN n18_CDNS_6738713766021 $T=105235 -19290 1 90 $X=104885 $Y=-19950
X487 GND 761 SAEN n18_CDNS_6738713766021 $T=109695 -19290 1 90 $X=109345 $Y=-19950
X488 INVB0 356 B0 343 ADD7 GND ICV_1 $T=42625 -9720 0 90 $X=41835 $Y=-10380
X489 INVB0 357 B0 344 ADD6 GND ICV_1 $T=42625 -3680 0 90 $X=41835 $Y=-4340
X490 INVB0 358 B0 345 ADD5 GND ICV_1 $T=42625 2360 0 90 $X=41835 $Y=1700
X491 INVB0 359 B0 346 ADD4 GND ICV_1 $T=42625 8400 0 90 $X=41835 $Y=7740
X492 INVB0 360 B0 347 ADD3 GND ICV_1 $T=42625 14440 0 90 $X=41835 $Y=13780
X493 INVB0 361 B0 348 ADD2 GND ICV_1 $T=42625 20480 0 90 $X=41835 $Y=19820
X494 INVB0 362 B0 349 ADD1 GND ICV_1 $T=42625 26520 0 90 $X=41835 $Y=25860
X495 INVB0 363 B0 350 ADD0 GND ICV_1 $T=42625 32560 0 90 $X=41835 $Y=31900
X496 INVB1 385 B1 372 ADD7 GND ICV_1 $T=47085 -9720 0 90 $X=46295 $Y=-10380
X497 INVB1 386 B1 373 ADD6 GND ICV_1 $T=47085 -3680 0 90 $X=46295 $Y=-4340
X498 INVB1 387 B1 374 ADD5 GND ICV_1 $T=47085 2360 0 90 $X=46295 $Y=1700
X499 INVB1 388 B1 375 ADD4 GND ICV_1 $T=47085 8400 0 90 $X=46295 $Y=7740
X500 INVB1 389 B1 376 ADD3 GND ICV_1 $T=47085 14440 0 90 $X=46295 $Y=13780
X501 INVB1 390 B1 377 ADD2 GND ICV_1 $T=47085 20480 0 90 $X=46295 $Y=19820
X502 INVB1 391 B1 378 ADD1 GND ICV_1 $T=47085 26520 0 90 $X=46295 $Y=25860
X503 INVB1 392 B1 379 ADD0 GND ICV_1 $T=47085 32560 0 90 $X=46295 $Y=31900
X504 INVB2 412 B2 399 ADD7 GND ICV_1 $T=51545 -9720 0 90 $X=50755 $Y=-10380
X505 INVB2 413 B2 400 ADD6 GND ICV_1 $T=51545 -3680 0 90 $X=50755 $Y=-4340
X506 INVB2 414 B2 401 ADD5 GND ICV_1 $T=51545 2360 0 90 $X=50755 $Y=1700
X507 INVB2 415 B2 402 ADD4 GND ICV_1 $T=51545 8400 0 90 $X=50755 $Y=7740
X508 INVB2 416 B2 403 ADD3 GND ICV_1 $T=51545 14440 0 90 $X=50755 $Y=13780
X509 INVB2 417 B2 404 ADD2 GND ICV_1 $T=51545 20480 0 90 $X=50755 $Y=19820
X510 INVB2 418 B2 405 ADD1 GND ICV_1 $T=51545 26520 0 90 $X=50755 $Y=25860
X511 INVB2 419 B2 406 ADD0 GND ICV_1 $T=51545 32560 0 90 $X=50755 $Y=31900
X512 INVB3 439 B3 426 ADD7 GND ICV_1 $T=56005 -9720 0 90 $X=55215 $Y=-10380
X513 INVB3 440 B3 427 ADD6 GND ICV_1 $T=56005 -3680 0 90 $X=55215 $Y=-4340
X514 INVB3 441 B3 428 ADD5 GND ICV_1 $T=56005 2360 0 90 $X=55215 $Y=1700
X515 INVB3 442 B3 429 ADD4 GND ICV_1 $T=56005 8400 0 90 $X=55215 $Y=7740
X516 INVB3 443 B3 430 ADD3 GND ICV_1 $T=56005 14440 0 90 $X=55215 $Y=13780
X517 INVB3 444 B3 431 ADD2 GND ICV_1 $T=56005 20480 0 90 $X=55215 $Y=19820
X518 INVB3 445 B3 432 ADD1 GND ICV_1 $T=56005 26520 0 90 $X=55215 $Y=25860
X519 INVB3 446 B3 433 ADD0 GND ICV_1 $T=56005 32560 0 90 $X=55215 $Y=31900
X520 INVB4 466 B4 453 ADD7 GND ICV_1 $T=60465 -9720 0 90 $X=59675 $Y=-10380
X521 INVB4 467 B4 454 ADD6 GND ICV_1 $T=60465 -3680 0 90 $X=59675 $Y=-4340
X522 INVB4 468 B4 455 ADD5 GND ICV_1 $T=60465 2360 0 90 $X=59675 $Y=1700
X523 INVB4 469 B4 456 ADD4 GND ICV_1 $T=60465 8400 0 90 $X=59675 $Y=7740
X524 INVB4 470 B4 457 ADD3 GND ICV_1 $T=60465 14440 0 90 $X=59675 $Y=13780
X525 INVB4 471 B4 458 ADD2 GND ICV_1 $T=60465 20480 0 90 $X=59675 $Y=19820
X526 INVB4 472 B4 459 ADD1 GND ICV_1 $T=60465 26520 0 90 $X=59675 $Y=25860
X527 INVB4 473 B4 460 ADD0 GND ICV_1 $T=60465 32560 0 90 $X=59675 $Y=31900
X528 INVB5 493 B5 482 ADD7 GND ICV_1 $T=64925 -9720 0 90 $X=64135 $Y=-10380
X529 INVB5 494 B5 483 ADD6 GND ICV_1 $T=64925 -3680 0 90 $X=64135 $Y=-4340
X530 INVB5 495 B5 484 ADD5 GND ICV_1 $T=64925 2360 0 90 $X=64135 $Y=1700
X531 INVB5 496 B5 485 ADD4 GND ICV_1 $T=64925 8400 0 90 $X=64135 $Y=7740
X532 INVB5 497 B5 486 ADD3 GND ICV_1 $T=64925 14440 0 90 $X=64135 $Y=13780
X533 INVB5 498 B5 487 ADD2 GND ICV_1 $T=64925 20480 0 90 $X=64135 $Y=19820
X534 INVB5 499 B5 488 ADD1 GND ICV_1 $T=64925 26520 0 90 $X=64135 $Y=25860
X535 INVB5 500 B5 489 ADD0 GND ICV_1 $T=64925 32560 0 90 $X=64135 $Y=31900
X536 INVB6 520 B6 509 ADD7 GND ICV_1 $T=69385 -9720 0 90 $X=68595 $Y=-10380
X537 INVB6 521 B6 510 ADD6 GND ICV_1 $T=69385 -3680 0 90 $X=68595 $Y=-4340
X538 INVB6 522 B6 511 ADD5 GND ICV_1 $T=69385 2360 0 90 $X=68595 $Y=1700
X539 INVB6 523 B6 512 ADD4 GND ICV_1 $T=69385 8400 0 90 $X=68595 $Y=7740
X540 INVB6 524 B6 513 ADD3 GND ICV_1 $T=69385 14440 0 90 $X=68595 $Y=13780
X541 INVB6 525 B6 514 ADD2 GND ICV_1 $T=69385 20480 0 90 $X=68595 $Y=19820
X542 INVB6 526 B6 515 ADD1 GND ICV_1 $T=69385 26520 0 90 $X=68595 $Y=25860
X543 INVB6 527 B6 516 ADD0 GND ICV_1 $T=69385 32560 0 90 $X=68595 $Y=31900
X544 INVB7 547 B7 536 ADD7 GND ICV_1 $T=73845 -9720 0 90 $X=73055 $Y=-10380
X545 INVB7 548 B7 537 ADD6 GND ICV_1 $T=73845 -3680 0 90 $X=73055 $Y=-4340
X546 INVB7 549 B7 538 ADD5 GND ICV_1 $T=73845 2360 0 90 $X=73055 $Y=1700
X547 INVB7 550 B7 539 ADD4 GND ICV_1 $T=73845 8400 0 90 $X=73055 $Y=7740
X548 INVB7 551 B7 540 ADD3 GND ICV_1 $T=73845 14440 0 90 $X=73055 $Y=13780
X549 INVB7 552 B7 541 ADD2 GND ICV_1 $T=73845 20480 0 90 $X=73055 $Y=19820
X550 INVB7 553 B7 542 ADD1 GND ICV_1 $T=73845 26520 0 90 $X=73055 $Y=25860
X551 INVB7 554 B7 543 ADD0 GND ICV_1 $T=73845 32560 0 90 $X=73055 $Y=31900
X552 INVB8 574 B8 563 ADD7 GND ICV_1 $T=78305 -9720 0 90 $X=77515 $Y=-10380
X553 INVB8 575 B8 564 ADD6 GND ICV_1 $T=78305 -3680 0 90 $X=77515 $Y=-4340
X554 INVB8 576 B8 565 ADD5 GND ICV_1 $T=78305 2360 0 90 $X=77515 $Y=1700
X555 INVB8 577 B8 566 ADD4 GND ICV_1 $T=78305 8400 0 90 $X=77515 $Y=7740
X556 INVB8 578 B8 567 ADD3 GND ICV_1 $T=78305 14440 0 90 $X=77515 $Y=13780
X557 INVB8 579 B8 568 ADD2 GND ICV_1 $T=78305 20480 0 90 $X=77515 $Y=19820
X558 INVB8 580 B8 569 ADD1 GND ICV_1 $T=78305 26520 0 90 $X=77515 $Y=25860
X559 INVB8 581 B8 570 ADD0 GND ICV_1 $T=78305 32560 0 90 $X=77515 $Y=31900
X560 INVB9 601 B9 590 ADD7 GND ICV_1 $T=82765 -9720 0 90 $X=81975 $Y=-10380
X561 INVB9 602 B9 591 ADD6 GND ICV_1 $T=82765 -3680 0 90 $X=81975 $Y=-4340
X562 INVB9 603 B9 592 ADD5 GND ICV_1 $T=82765 2360 0 90 $X=81975 $Y=1700
X563 INVB9 604 B9 593 ADD4 GND ICV_1 $T=82765 8400 0 90 $X=81975 $Y=7740
X564 INVB9 605 B9 594 ADD3 GND ICV_1 $T=82765 14440 0 90 $X=81975 $Y=13780
X565 INVB9 606 B9 595 ADD2 GND ICV_1 $T=82765 20480 0 90 $X=81975 $Y=19820
X566 INVB9 607 B9 596 ADD1 GND ICV_1 $T=82765 26520 0 90 $X=81975 $Y=25860
X567 INVB9 608 B9 597 ADD0 GND ICV_1 $T=82765 32560 0 90 $X=81975 $Y=31900
X568 INVB10 630 B10 617 ADD7 GND ICV_1 $T=87225 -9720 0 90 $X=86435 $Y=-10380
X569 INVB10 631 B10 618 ADD6 GND ICV_1 $T=87225 -3680 0 90 $X=86435 $Y=-4340
X570 INVB10 632 B10 619 ADD5 GND ICV_1 $T=87225 2360 0 90 $X=86435 $Y=1700
X571 INVB10 633 B10 620 ADD4 GND ICV_1 $T=87225 8400 0 90 $X=86435 $Y=7740
X572 INVB10 634 B10 621 ADD3 GND ICV_1 $T=87225 14440 0 90 $X=86435 $Y=13780
X573 INVB10 635 B10 622 ADD2 GND ICV_1 $T=87225 20480 0 90 $X=86435 $Y=19820
X574 INVB10 636 B10 623 ADD1 GND ICV_1 $T=87225 26520 0 90 $X=86435 $Y=25860
X575 INVB10 637 B10 624 ADD0 GND ICV_1 $T=87225 32560 0 90 $X=86435 $Y=31900
X576 INVB11 657 B11 644 ADD7 GND ICV_1 $T=91685 -9720 0 90 $X=90895 $Y=-10380
X577 INVB11 658 B11 645 ADD6 GND ICV_1 $T=91685 -3680 0 90 $X=90895 $Y=-4340
X578 INVB11 659 B11 646 ADD5 GND ICV_1 $T=91685 2360 0 90 $X=90895 $Y=1700
X579 INVB11 660 B11 647 ADD4 GND ICV_1 $T=91685 8400 0 90 $X=90895 $Y=7740
X580 INVB11 661 B11 648 ADD3 GND ICV_1 $T=91685 14440 0 90 $X=90895 $Y=13780
X581 INVB11 662 B11 649 ADD2 GND ICV_1 $T=91685 20480 0 90 $X=90895 $Y=19820
X582 INVB11 663 B11 650 ADD1 GND ICV_1 $T=91685 26520 0 90 $X=90895 $Y=25860
X583 INVB11 664 B11 651 ADD0 GND ICV_1 $T=91685 32560 0 90 $X=90895 $Y=31900
X584 INVB12 686 B12 673 ADD7 GND ICV_1 $T=96145 -9720 0 90 $X=95355 $Y=-10380
X585 INVB12 687 B12 674 ADD6 GND ICV_1 $T=96145 -3680 0 90 $X=95355 $Y=-4340
X586 INVB12 688 B12 675 ADD5 GND ICV_1 $T=96145 2360 0 90 $X=95355 $Y=1700
X587 INVB12 689 B12 676 ADD4 GND ICV_1 $T=96145 8400 0 90 $X=95355 $Y=7740
X588 INVB12 690 B12 677 ADD3 GND ICV_1 $T=96145 14440 0 90 $X=95355 $Y=13780
X589 INVB12 691 B12 678 ADD2 GND ICV_1 $T=96145 20480 0 90 $X=95355 $Y=19820
X590 INVB12 692 B12 679 ADD1 GND ICV_1 $T=96145 26520 0 90 $X=95355 $Y=25860
X591 INVB12 693 B12 680 ADD0 GND ICV_1 $T=96145 32560 0 90 $X=95355 $Y=31900
X592 INVB13 711 B13 700 ADD7 GND ICV_1 $T=100605 -9720 0 90 $X=99815 $Y=-10380
X593 INVB13 712 B13 701 ADD6 GND ICV_1 $T=100605 -3680 0 90 $X=99815 $Y=-4340
X594 INVB13 713 B13 702 ADD5 GND ICV_1 $T=100605 2360 0 90 $X=99815 $Y=1700
X595 INVB13 714 B13 703 ADD4 GND ICV_1 $T=100605 8400 0 90 $X=99815 $Y=7740
X596 INVB13 715 B13 704 ADD3 GND ICV_1 $T=100605 14440 0 90 $X=99815 $Y=13780
X597 INVB13 716 B13 705 ADD2 GND ICV_1 $T=100605 20480 0 90 $X=99815 $Y=19820
X598 INVB13 717 B13 706 ADD1 GND ICV_1 $T=100605 26520 0 90 $X=99815 $Y=25860
X599 INVB13 718 B13 707 ADD0 GND ICV_1 $T=100605 32560 0 90 $X=99815 $Y=31900
X600 INVB14 740 B14 727 ADD7 GND ICV_1 $T=105065 -9720 0 90 $X=104275 $Y=-10380
X601 INVB14 741 B14 728 ADD6 GND ICV_1 $T=105065 -3680 0 90 $X=104275 $Y=-4340
X602 INVB14 742 B14 729 ADD5 GND ICV_1 $T=105065 2360 0 90 $X=104275 $Y=1700
X603 INVB14 743 B14 730 ADD4 GND ICV_1 $T=105065 8400 0 90 $X=104275 $Y=7740
X604 INVB14 744 B14 731 ADD3 GND ICV_1 $T=105065 14440 0 90 $X=104275 $Y=13780
X605 INVB14 745 B14 732 ADD2 GND ICV_1 $T=105065 20480 0 90 $X=104275 $Y=19820
X606 INVB14 746 B14 733 ADD1 GND ICV_1 $T=105065 26520 0 90 $X=104275 $Y=25860
X607 INVB14 747 B14 734 ADD0 GND ICV_1 $T=105065 32560 0 90 $X=104275 $Y=31900
X608 INVB15 763 B15 752 ADD7 GND ICV_1 $T=109525 -9720 0 90 $X=108735 $Y=-10380
X609 INVB15 764 B15 753 ADD6 GND ICV_1 $T=109525 -3680 0 90 $X=108735 $Y=-4340
X610 INVB15 765 B15 754 ADD5 GND ICV_1 $T=109525 2360 0 90 $X=108735 $Y=1700
X611 INVB15 766 B15 755 ADD4 GND ICV_1 $T=109525 8400 0 90 $X=108735 $Y=7740
X612 INVB15 767 B15 756 ADD3 GND ICV_1 $T=109525 14440 0 90 $X=108735 $Y=13780
X613 INVB15 768 B15 757 ADD2 GND ICV_1 $T=109525 20480 0 90 $X=108735 $Y=19820
X614 INVB15 769 B15 758 ADD1 GND ICV_1 $T=109525 26520 0 90 $X=108735 $Y=25860
X615 INVB15 770 B15 759 ADD0 GND ICV_1 $T=109525 32560 0 90 $X=108735 $Y=31900
X616 GND 340 B0 INVB0 367 368 B1 INVB1 394 94 MODE 98 99 102 ICV_3 $T=42135 -32390 0 0 $X=41475 $Y=-33520
X617 GND 395 B2 INVB2 421 422 B3 INVB3 448 103 MODE 106 107 110 ICV_3 $T=51055 -32390 0 0 $X=50395 $Y=-33520
X618 GND 451 B4 INVB4 475 478 B5 INVB5 502 111 MODE 114 115 118 ICV_3 $T=59975 -32390 0 0 $X=59315 $Y=-33520
X619 GND 505 B6 INVB6 529 534 B7 INVB7 558 119 MODE 122 124 127 ICV_3 $T=68895 -32390 0 0 $X=68235 $Y=-33520
X620 GND 561 B8 INVB8 585 588 B9 INVB9 612 128 MODE 131 132 135 ICV_3 $T=77815 -32390 0 0 $X=77155 $Y=-33520
X621 GND 615 B10 INVB10 641 642 B11 INVB11 666 136 MODE 139 140 143 ICV_3 $T=86735 -32390 0 0 $X=86075 $Y=-33520
X622 GND 669 B12 INVB12 695 696 B13 INVB13 722 144 MODE 147 148 151 ICV_3 $T=95655 -32390 0 0 $X=94995 $Y=-33520
X623 GND 723 B14 INVB14 749 750 B15 INVB15 772 152 MODE 155 156 159 ICV_3 $T=104575 -32390 0 0 $X=103915 $Y=-33520
X624 VDD VDD 28 A2 p18_CDNS_673871376605 $T=-16580 -1400 1 270 $X=-18150 $Y=-2490
X625 VDD VDD 30 A1 p18_CDNS_673871376605 $T=-16580 620 1 270 $X=-18150 $Y=-470
X626 VDD VDD 29 A0 p18_CDNS_673871376605 $T=-16580 2640 1 270 $X=-18150 $Y=1550
X627 VDD VDD 1 194 p18_CDNS_673871376605 $T=-6135 -9600 1 270 $X=-7705 $Y=-10690
X628 VDD VDD 6 195 p18_CDNS_673871376605 $T=-6135 -4960 1 270 $X=-7705 $Y=-6050
X629 VDD VDD 5 196 p18_CDNS_673871376605 $T=-6135 -320 1 270 $X=-7705 $Y=-1410
X630 VDD VDD 7 197 p18_CDNS_673871376605 $T=-6135 4320 1 270 $X=-7705 $Y=3230
X631 VDD VDD 8 198 p18_CDNS_673871376605 $T=-6135 8960 1 270 $X=-7705 $Y=7870
X632 VDD VDD 2 201 p18_CDNS_673871376605 $T=-6135 22880 1 270 $X=-7705 $Y=21790
X633 VDD VDD 296 285 p18_CDNS_673871376605 $T=20495 47490 0 0 $X=19585 $Y=47060
X634 VDD VDD 52 50 p18_CDNS_673871376605 $T=25135 -26350 1 0 $X=24225 $Y=-27920
X635 VDD VDD 53 306 p18_CDNS_673871376605 $T=25135 47490 0 0 $X=24225 $Y=47060
X636 VDD VDD 55 VDD p18_CDNS_673871376605 $T=27155 47490 0 0 $X=26245 $Y=47060
X637 VDD VDD 64 MODE p18_CDNS_673871376605 $T=29175 -26350 1 0 $X=28265 $Y=-27920
X638 VDD VDD 65 MODE p18_CDNS_673871376605 $T=29175 47490 0 0 $X=28265 $Y=47060
X639 VDD VDD 327 326 p18_CDNS_673871376605 $T=34495 -28710 0 0 $X=33585 $Y=-29140
X640 VDD B0 INVB0 B1 INVB1 PCEN ICV_5 $T=42175 39870 0 0 $X=41265 $Y=39440
X641 VDD B2 INVB2 B3 INVB3 PCEN ICV_5 $T=51095 39870 0 0 $X=50185 $Y=39440
X642 VDD B4 INVB4 B5 INVB5 PCEN ICV_5 $T=60015 39870 0 0 $X=59105 $Y=39440
X643 VDD B6 INVB6 B7 INVB7 PCEN ICV_5 $T=68935 39870 0 0 $X=68025 $Y=39440
X644 VDD B8 INVB8 B9 INVB9 PCEN ICV_5 $T=77855 39870 0 0 $X=76945 $Y=39440
X645 VDD B10 INVB10 B11 INVB11 PCEN ICV_5 $T=86775 39870 0 0 $X=85865 $Y=39440
X646 VDD B12 INVB12 B13 INVB13 PCEN ICV_5 $T=95695 39870 0 0 $X=94785 $Y=39440
X647 VDD B14 INVB14 B15 INVB15 PCEN ICV_5 $T=104615 39870 0 0 $X=103705 $Y=39440
X648 VDD 384 10 355 9 GND 393 364 ICV_8 $T=42315 -22610 1 180 $X=41225 $Y=-23740
X649 VDD 438 12 411 11 GND 447 420 ICV_8 $T=51235 -22610 1 180 $X=50145 $Y=-23740
X650 VDD 492 14 465 13 GND 501 474 ICV_8 $T=60155 -22610 1 180 $X=59065 $Y=-23740
X651 VDD 546 16 519 15 GND 555 528 ICV_8 $T=69075 -22610 1 180 $X=67985 $Y=-23740
X652 VDD 600 18 573 17 GND 611 584 ICV_8 $T=77995 -22610 1 180 $X=76905 $Y=-23740
X653 VDD 656 20 629 19 GND 665 638 ICV_8 $T=86915 -22610 1 180 $X=85825 $Y=-23740
X654 VDD 710 22 685 21 GND 721 694 ICV_8 $T=95835 -22610 1 180 $X=94745 $Y=-23740
X655 VDD 762 24 739 23 GND 771 748 ICV_8 $T=104755 -22610 1 180 $X=103665 $Y=-23740
X656 GND VDD 343 356 372 385 399 412 426 439 453 466 482 493 509 520 536 547 563 574
+ 590 601 617 630 644 657 673 686 700 711 727 740 752 763
+ ICV_15 $T=42135 -8090 0 0 $X=40615 $Y=-8440
X657 GND VDD 344 357 373 386 400 413 427 440 454 467 483 494 510 521 537 548 564 575
+ 591 602 618 631 645 658 674 687 701 712 728 741 753 764
+ ICV_15 $T=42135 -2050 0 0 $X=40615 $Y=-2400
X658 GND VDD 345 358 374 387 401 414 428 441 455 468 484 495 511 522 538 549 565 576
+ 592 603 619 632 646 659 675 688 702 713 729 742 754 765
+ ICV_15 $T=42135 3990 0 0 $X=40615 $Y=3640
X659 GND VDD 346 359 375 388 402 415 429 442 456 469 485 496 512 523 539 550 566 577
+ 593 604 620 633 647 660 676 689 703 714 730 743 755 766
+ ICV_15 $T=42135 10030 0 0 $X=40615 $Y=9680
X660 GND VDD 347 360 376 389 403 416 430 443 457 470 486 497 513 524 540 551 567 578
+ 594 605 621 634 648 661 677 690 704 715 731 744 756 767
+ ICV_15 $T=42135 16070 0 0 $X=40615 $Y=15720
X661 GND VDD 348 361 377 390 404 417 431 444 458 471 487 498 514 525 541 552 568 579
+ 595 606 622 635 649 662 678 691 705 716 732 745 757 768
+ ICV_15 $T=42135 22110 0 0 $X=40615 $Y=21760
X662 GND VDD 349 362 378 391 405 418 432 445 459 472 488 499 515 526 542 553 569 580
+ 596 607 623 636 650 663 679 692 706 717 733 746 758 769
+ ICV_15 $T=42135 28150 0 0 $X=40615 $Y=27800
X663 GND VDD 350 363 379 392 406 419 433 446 460 473 489 500 516 527 543 554 570 581
+ 597 608 624 637 651 664 680 693 707 718 734 747 759 770
+ ICV_15 $T=42135 34190 0 0 $X=40615 $Y=33840
X664 GND 328 327 n18_CDNS_6738713766013 $T=36475 -34410 0 0 $X=35815 $Y=-35540
X665 GND CLKREG 328 n18_CDNS_6738713766013 $T=38415 -34410 0 0 $X=37755 $Y=-35540
X666 VDD 328 327 p18_CDNS_6738713766014 $T=36475 -31790 0 0 $X=35565 $Y=-32220
X667 VDD CLKREG 328 p18_CDNS_6738713766014 $T=38415 -31790 0 0 $X=37505 $Y=-32220
X668 GND 40 74 MODE n18_CDNS_6738713766011 $T=31155 -20650 1 0 $X=30495 $Y=-21440
X669 GND ADD7 85 MODE n18_CDNS_6738713766011 $T=35035 -19170 0 0 $X=34375 $Y=-20300
X670 GND ADD6 86 MODE n18_CDNS_6738713766011 $T=35035 -5410 1 0 $X=34375 $Y=-6200
X671 GND ADD5 87 MODE n18_CDNS_6738713766011 $T=35035 -3930 0 0 $X=34375 $Y=-5060
X672 GND ADD4 88 MODE n18_CDNS_6738713766011 $T=35035 9830 1 0 $X=34375 $Y=9040
X673 GND ADD3 89 MODE n18_CDNS_6738713766011 $T=35035 11310 0 0 $X=34375 $Y=10180
X674 GND ADD2 90 MODE n18_CDNS_6738713766011 $T=35035 25070 1 0 $X=34375 $Y=24280
X675 GND ADD1 91 MODE n18_CDNS_6738713766011 $T=35035 26550 0 0 $X=34375 $Y=25420
X676 GND ADD0 92 MODE n18_CDNS_6738713766011 $T=35035 40310 1 0 $X=34375 $Y=39520
X677 GND GND 85 66 n18_CDNS_6738713766011 $T=37695 -19170 0 0 $X=37035 $Y=-20300
X678 GND GND 86 67 n18_CDNS_6738713766011 $T=37695 -5410 1 0 $X=37035 $Y=-6200
X679 GND GND 87 68 n18_CDNS_6738713766011 $T=37695 -3930 0 0 $X=37035 $Y=-5060
X680 GND GND 88 69 n18_CDNS_6738713766011 $T=37695 9830 1 0 $X=37035 $Y=9040
X681 GND GND 89 70 n18_CDNS_6738713766011 $T=37695 11310 0 0 $X=37035 $Y=10180
X682 GND GND 90 71 n18_CDNS_6738713766011 $T=37695 25070 1 0 $X=37035 $Y=24280
X683 GND GND 91 72 n18_CDNS_6738713766011 $T=37695 26550 0 0 $X=37035 $Y=25420
X684 GND 329 40 n18_CDNS_673871376608 $T=36475 -20650 1 0 $X=35815 $Y=-21880
X685 GND 204 214 203 ICV_16 $T=1055 41790 0 0 $X=395 $Y=40660
X686 GND 257 268 247 ICV_16 $T=13795 -19170 0 0 $X=13135 $Y=-20300
X687 GND 50 267 256 ICV_16 $T=14635 41790 0 0 $X=13975 $Y=40660
X688 GND 307 324 297 ICV_16 $T=25935 -34410 0 0 $X=25275 $Y=-35540
X689 GND 330 PCEN 41 ICV_16 $T=36475 41790 0 0 $X=35815 $Y=40660
X690 VDD 324 307 p18_CDNS_673871376609 $T=27875 -30030 0 0 $X=26965 $Y=-30460
X691 VDD 267 285 50 ICV_17 $T=16575 46170 0 0 $X=15665 $Y=45740
X692 VDD 329 SAEN 40 ICV_17 $T=36475 -25030 1 0 $X=35565 $Y=-27920
X693 VDD 330 PCEN 41 ICV_17 $T=36475 46170 0 0 $X=35565 $Y=45740
X694 VDD MODE 832 p18_CDNS_6738713766010 $T=31155 -25910 1 0 $X=30245 $Y=-27920
X695 VDD 41 MODE 53 ICV_18 $T=31155 47050 0 0 $X=30245 $Y=46620
X696 VDD ADD7 MODE 56 ICV_18 $T=35035 -13910 0 0 $X=34125 $Y=-14340
X697 VDD ADD6 MODE 57 ICV_18 $T=35035 -10670 1 0 $X=34125 $Y=-12680
X698 VDD ADD5 MODE 58 ICV_18 $T=35035 1330 0 0 $X=34125 $Y=900
X699 VDD ADD4 MODE 59 ICV_18 $T=35035 4570 1 0 $X=34125 $Y=2560
X700 VDD ADD3 MODE 60 ICV_18 $T=35035 16570 0 0 $X=34125 $Y=16140
X701 VDD ADD2 MODE 61 ICV_18 $T=35035 19810 1 0 $X=34125 $Y=17800
X702 VDD ADD1 MODE 62 ICV_18 $T=35035 31810 0 0 $X=34125 $Y=31380
X703 VDD ADD0 MODE 63 ICV_18 $T=35035 35050 1 0 $X=34125 $Y=33040
X704 GND 205 41 n18_CDNS_673871376606 $T=2035 -19070 0 0 $X=1335 $Y=-20300
X705 GND 42 205 n18_CDNS_673871376606 $T=4055 -19070 0 0 $X=3355 $Y=-20300
X706 GND 276 268 n18_CDNS_673871376606 $T=17715 -19070 0 0 $X=17015 $Y=-20300
X707 GND 283 275 n18_CDNS_673871376606 $T=17715 40210 1 0 $X=17015 $Y=39640
X708 GND 296 285 n18_CDNS_673871376606 $T=20495 41890 0 0 $X=19795 $Y=40660
X709 GND 298 287 n18_CDNS_673871376606 $T=22355 -19070 0 0 $X=21655 $Y=-20300
X710 GND 305 294 n18_CDNS_673871376606 $T=22355 40210 1 0 $X=21655 $Y=39640
X711 GND 52 50 n18_CDNS_673871376606 $T=25135 -20750 1 0 $X=24435 $Y=-21320
X712 GND 53 306 n18_CDNS_673871376606 $T=25135 41890 0 0 $X=24435 $Y=40660
X713 GND 54 GND n18_CDNS_673871376606 $T=27155 -20750 1 0 $X=26455 $Y=-21320
X714 GND 55 VDD n18_CDNS_673871376606 $T=27155 41890 0 0 $X=26455 $Y=40660
X715 GND 64 MODE n18_CDNS_673871376606 $T=29175 -20750 1 0 $X=28475 $Y=-21320
X716 GND 65 MODE n18_CDNS_673871376606 $T=29175 41890 0 0 $X=28475 $Y=40660
X717 GND 325 324 n18_CDNS_673871376606 $T=29855 -34310 0 0 $X=29155 $Y=-35540
X718 GND 73 2 n18_CDNS_673871376606 $T=31035 40210 1 0 $X=30335 $Y=39640
X719 GND 77 MODE n18_CDNS_673871376606 $T=33055 -19070 0 0 $X=32355 $Y=-20300
X720 GND 84 MODE n18_CDNS_673871376606 $T=33055 40210 1 0 $X=32355 $Y=39640
X721 GND 327 326 n18_CDNS_673871376606 $T=34495 -34310 0 0 $X=33795 $Y=-35540
X722 GND 287 42 809 n18_CDNS_673871376600 $T=20125 -19170 0 0 $X=19805 $Y=-20300
X723 GND 288 43 810 n18_CDNS_673871376600 $T=20125 -5410 1 0 $X=19805 $Y=-6200
X724 GND 289 44 811 n18_CDNS_673871376600 $T=20125 -3930 0 0 $X=19805 $Y=-5060
X725 GND 290 45 812 n18_CDNS_673871376600 $T=20125 9830 1 0 $X=19805 $Y=9040
X726 GND 291 46 813 n18_CDNS_673871376600 $T=20125 11310 0 0 $X=19805 $Y=10180
X727 GND 292 47 814 n18_CDNS_673871376600 $T=20125 25070 1 0 $X=19805 $Y=24280
X728 GND 293 48 815 n18_CDNS_673871376600 $T=20125 26550 0 0 $X=19805 $Y=25420
X729 GND 309 299 816 n18_CDNS_673871376600 $T=24765 -5410 1 0 $X=24445 $Y=-6200
X730 GND 310 300 817 n18_CDNS_673871376600 $T=24765 -3930 0 0 $X=24445 $Y=-5060
X731 GND 311 301 818 n18_CDNS_673871376600 $T=24765 9830 1 0 $X=24445 $Y=9040
X732 GND 312 302 819 n18_CDNS_673871376600 $T=24765 11310 0 0 $X=24445 $Y=10180
X733 GND 313 303 820 n18_CDNS_673871376600 $T=24765 25070 1 0 $X=24445 $Y=24280
X734 GND 314 304 821 n18_CDNS_673871376600 $T=24765 26550 0 0 $X=24445 $Y=25420
X735 GND 326 325 822 n18_CDNS_673871376600 $T=32265 -34410 0 0 $X=31945 $Y=-35540
X736 GND 276 809 n18_CDNS_673871376601 $T=19695 -19170 0 0 $X=19035 $Y=-20300
X737 GND 277 810 n18_CDNS_673871376601 $T=19695 -5410 1 0 $X=19035 $Y=-6200
X738 GND 278 811 n18_CDNS_673871376601 $T=19695 -3930 0 0 $X=19035 $Y=-5060
X739 GND 279 812 n18_CDNS_673871376601 $T=19695 9830 1 0 $X=19035 $Y=9040
X740 GND 280 813 n18_CDNS_673871376601 $T=19695 11310 0 0 $X=19035 $Y=10180
X741 GND 281 814 n18_CDNS_673871376601 $T=19695 25070 1 0 $X=19035 $Y=24280
X742 GND 282 815 n18_CDNS_673871376601 $T=19695 26550 0 0 $X=19035 $Y=25420
X743 GND 283 773 n18_CDNS_673871376601 $T=19695 40310 1 0 $X=19035 $Y=39520
X744 GND 1 775 n18_CDNS_673871376601 $T=24335 -19170 0 0 $X=23675 $Y=-20300
X745 GND 6 816 n18_CDNS_673871376601 $T=24335 -5410 1 0 $X=23675 $Y=-6200
X746 GND 5 817 n18_CDNS_673871376601 $T=24335 -3930 0 0 $X=23675 $Y=-5060
X747 GND 7 818 n18_CDNS_673871376601 $T=24335 9830 1 0 $X=23675 $Y=9040
X748 GND 8 819 n18_CDNS_673871376601 $T=24335 11310 0 0 $X=23675 $Y=10180
X749 GND 4 820 n18_CDNS_673871376601 $T=24335 25070 1 0 $X=23675 $Y=24280
X750 GND 3 821 n18_CDNS_673871376601 $T=24335 26550 0 0 $X=23675 $Y=25420
X751 GND 2 776 n18_CDNS_673871376601 $T=24335 40310 1 0 $X=23675 $Y=39520
X752 GND 76 822 n18_CDNS_673871376601 $T=31835 -34410 0 0 $X=31175 $Y=-35540
X753 VDD 194 CLK p18_CDNS_673871376607 $T=-5695 -6940 1 270 $X=-7705 $Y=-8030
X754 VDD 195 CLK p18_CDNS_673871376607 $T=-5695 -2300 1 270 $X=-7705 $Y=-3390
X755 VDD 196 CLK p18_CDNS_673871376607 $T=-5695 2340 1 270 $X=-7705 $Y=1250
X756 VDD 197 CLK p18_CDNS_673871376607 $T=-5695 6980 1 270 $X=-7705 $Y=5890
X757 VDD 198 CLK p18_CDNS_673871376607 $T=-5695 11620 1 270 $X=-7705 $Y=10530
X758 VDD 199 CLK p18_CDNS_673871376607 $T=-5695 16260 1 270 $X=-7705 $Y=15170
X759 VDD 306 CLK p18_CDNS_673871376607 $T=22475 47050 0 0 $X=21565 $Y=46620
X760 VDD 326 76 p18_CDNS_673871376607 $T=31835 -29150 0 0 $X=30925 $Y=-29580
X761 GND 278 277 270 269 ICV_19 $T=17715 -5510 1 0 $X=17015 $Y=-6080
X762 GND 280 279 272 271 ICV_19 $T=17715 9730 1 0 $X=17015 $Y=9160
X763 GND 282 281 274 273 ICV_19 $T=17715 24970 1 0 $X=17015 $Y=24400
X764 GND 300 299 289 288 ICV_19 $T=22355 -5510 1 0 $X=21655 $Y=-6080
X765 GND 302 301 291 290 ICV_19 $T=22355 9730 1 0 $X=21655 $Y=9160
X766 GND 304 303 293 292 ICV_19 $T=22355 24970 1 0 $X=21655 $Y=24400
X767 GND 207 206 44 43 41 41 207 206 ICV_20 $T=2035 -5510 1 0 $X=1335 $Y=-6080
X768 GND 209 208 46 45 41 41 209 208 ICV_20 $T=2035 9730 1 0 $X=1335 $Y=9160
X769 GND 211 210 48 47 41 41 211 210 ICV_20 $T=2035 24970 1 0 $X=1335 $Y=24400
X770 GND 318 317 58 57 310 309 318 317 ICV_20 $T=26995 -5510 1 0 $X=26295 $Y=-6080
X771 GND 320 319 60 59 312 311 320 319 ICV_20 $T=26995 9730 1 0 $X=26295 $Y=9160
X772 GND 322 321 62 61 314 313 322 321 ICV_20 $T=26995 24970 1 0 $X=26295 $Y=24400
X773 GND 68 67 79 78 5 6 MODE MODE ICV_20 $T=31035 -5510 1 0 $X=30335 $Y=-6080
X774 GND 70 69 81 80 8 7 MODE MODE ICV_20 $T=31035 9730 1 0 $X=30335 $Y=9160
X775 GND 72 71 83 82 3 4 MODE MODE ICV_20 $T=31035 24970 1 0 $X=30335 $Y=24400
X776 VDD 276 277 268 269 ICV_21 $T=17715 -13470 0 0 $X=16805 $Y=-13900
X777 VDD 278 279 270 271 ICV_21 $T=17715 1770 0 0 $X=16805 $Y=1340
X778 VDD 280 281 272 273 ICV_21 $T=17715 17010 0 0 $X=16805 $Y=16580
X779 VDD 282 283 274 275 ICV_21 $T=17715 32250 0 0 $X=16805 $Y=31820
X780 VDD 298 299 287 288 ICV_21 $T=22355 -13470 0 0 $X=21445 $Y=-13900
X781 VDD 300 301 289 290 ICV_21 $T=22355 1770 0 0 $X=21445 $Y=1340
X782 VDD 302 303 291 292 ICV_21 $T=22355 17010 0 0 $X=21445 $Y=16580
X783 VDD 304 305 293 294 ICV_21 $T=22355 32250 0 0 $X=21445 $Y=31820
X784 VDD 205 206 42 43 41 41 205 206 ICV_22 $T=2035 -13470 0 0 $X=1125 $Y=-13900
X785 VDD 207 208 44 45 41 41 207 208 ICV_22 $T=2035 1770 0 0 $X=1125 $Y=1340
X786 VDD 209 210 46 47 41 41 209 210 ICV_22 $T=2035 17010 0 0 $X=1125 $Y=16580
X787 VDD 211 212 48 49 41 41 211 212 ICV_22 $T=2035 32250 0 0 $X=1125 $Y=31820
X788 VDD 316 317 56 57 308 309 316 317 ICV_22 $T=26995 -13470 0 0 $X=26085 $Y=-13900
X789 VDD 318 319 58 59 310 311 318 319 ICV_22 $T=26995 1770 0 0 $X=26085 $Y=1340
X790 VDD 320 321 60 61 312 313 320 321 ICV_22 $T=26995 17010 0 0 $X=26085 $Y=16580
X791 VDD 322 323 62 63 314 315 322 323 ICV_22 $T=26995 32250 0 0 $X=26085 $Y=31820
X792 VDD 66 67 77 78 1 6 MODE MODE ICV_22 $T=31035 -13470 0 0 $X=30125 $Y=-13900
X793 VDD 68 69 79 80 5 7 MODE MODE ICV_22 $T=31035 1770 0 0 $X=30125 $Y=1340
X794 VDD 70 71 81 82 8 4 MODE MODE ICV_22 $T=31035 17010 0 0 $X=30125 $Y=16580
X795 VDD 72 73 83 84 3 2 MODE MODE ICV_22 $T=31035 32250 0 0 $X=30125 $Y=31820
X796 VDD 287 288 276 277 ICV_23 $T=19695 -13910 0 0 $X=18785 $Y=-14340
X797 VDD 289 290 278 279 ICV_23 $T=19695 1330 0 0 $X=18785 $Y=900
X798 VDD 291 292 280 281 ICV_23 $T=19695 16570 0 0 $X=18785 $Y=16140
X799 VDD 293 294 282 283 ICV_23 $T=19695 31810 0 0 $X=18785 $Y=31380
X800 VDD 308 309 1 6 ICV_23 $T=24335 -13910 0 0 $X=23425 $Y=-14340
X801 VDD 310 311 5 7 ICV_23 $T=24335 1330 0 0 $X=23425 $Y=900
X802 VDD 312 313 8 4 ICV_23 $T=24335 16570 0 0 $X=23425 $Y=16140
X803 VDD 314 315 3 2 ICV_23 $T=24335 31810 0 0 $X=23425 $Y=31380
X804 GND 219 218 229 228 44 43 ICV_25 $T=6035 -5410 1 0 $X=5375 $Y=-6640
X805 GND 221 220 231 230 46 45 ICV_25 $T=6035 9830 1 0 $X=5375 $Y=8600
X806 GND 223 222 233 232 48 47 ICV_25 $T=6035 25070 1 0 $X=5375 $Y=23840
X807 GND 239 238 249 248 229 228 ICV_25 $T=9915 -5410 1 0 $X=9255 $Y=-6640
X808 GND 241 240 251 250 231 230 ICV_25 $T=9915 9830 1 0 $X=9255 $Y=8600
X809 GND 243 242 253 252 233 232 ICV_25 $T=9915 25070 1 0 $X=9255 $Y=23840
X810 GND 259 258 270 269 249 248 ICV_25 $T=13795 -5410 1 0 $X=13135 $Y=-6640
X811 GND 261 260 272 271 251 250 ICV_25 $T=13795 9830 1 0 $X=13135 $Y=8600
X812 GND 263 262 274 273 253 252 ICV_25 $T=13795 25070 1 0 $X=13135 $Y=23840
X813 VDD 257 268 258 269 247 248 ICV_26 $T=13795 -14790 0 0 $X=12885 $Y=-15220
X814 VDD 259 270 260 271 249 250 ICV_26 $T=13795 450 0 0 $X=12885 $Y=20
X815 VDD 261 272 262 273 251 252 ICV_26 $T=13795 15690 0 0 $X=12885 $Y=15260
X816 VDD 263 274 264 275 253 254 ICV_26 $T=13795 30930 0 0 $X=12885 $Y=30500
X817 GND 217 227 237 247 42 ICV_27 $T=6035 -19170 0 0 $X=5375 $Y=-20300
X818 GND 226 236 246 256 216 ICV_27 $T=6875 41790 0 0 $X=6215 $Y=40660
X819 GND 161 162 163 164 165 166 167 168 40 ICV_28 $T=-51665 -34410 0 0 $X=-52325 $Y=-35540
X820 GND 169 170 171 172 173 174 175 176 168 ICV_28 $T=-36145 -34410 0 0 $X=-36805 $Y=-35540
X821 GND 177 178 179 180 182 184 186 188 176 ICV_28 $T=-20625 -34410 0 0 $X=-21285 $Y=-35540
X822 GND 181 183 185 187 189 191 193 203 CLK ICV_28 $T=-14465 41790 0 0 $X=-15125 $Y=40660
X823 GND 190 192 202 76 213 215 225 235 188 ICV_28 $T=-5105 -34410 0 0 $X=-5765 $Y=-35540
X824 GND 245 255 265 266 284 286 295 297 235 ICV_28 $T=10415 -34410 0 0 $X=9755 $Y=-35540
X825 VDD 161 162 163 164 165 166 167 168 40 ICV_30 $T=-51665 -30030 0 0 $X=-52575 $Y=-30460
X826 VDD 169 170 171 172 173 174 175 176 168 ICV_30 $T=-36145 -30030 0 0 $X=-37055 $Y=-30460
X827 VDD 177 178 179 180 182 184 186 188 176 ICV_30 $T=-20625 -30030 0 0 $X=-21535 $Y=-30460
X828 VDD 181 183 185 187 189 191 193 203 CLK ICV_30 $T=-14465 46170 0 0 $X=-15375 $Y=45740
X829 VDD 190 192 202 76 213 215 225 235 188 ICV_30 $T=-5105 -30030 0 0 $X=-6015 $Y=-30460
X830 VDD 204 214 216 226 236 246 256 50 203 ICV_30 $T=1055 46170 0 0 $X=145 $Y=45740
X831 VDD 245 255 265 266 284 286 295 297 235 ICV_30 $T=10415 -30030 0 0 $X=9505 $Y=-30460
X832 VDD 217 218 227 228 237 238 247 248 42 43 ICV_31 $T=6035 -14790 0 0 $X=5125 $Y=-15220
X833 VDD 219 220 229 230 239 240 249 250 44 45 ICV_31 $T=6035 450 0 0 $X=5125 $Y=20
X834 VDD 221 222 231 232 241 242 251 252 46 47 ICV_31 $T=6035 15690 0 0 $X=5125 $Y=15260
X835 VDD 223 224 233 234 243 244 253 254 48 49 ICV_31 $T=6035 30930 0 0 $X=5125 $Y=30500
X836 GND 1 194 31 CLK ICV_32 $T=-535 -9600 1 270 $X=-1225 $Y=-10480
X837 GND 6 195 34 CLK ICV_32 $T=-535 -4960 1 270 $X=-1225 $Y=-5840
X838 GND 5 196 35 CLK ICV_32 $T=-535 -320 1 270 $X=-1225 $Y=-1200
X839 GND 7 197 36 CLK ICV_32 $T=-535 4320 1 270 $X=-1225 $Y=3440
X840 GND 8 198 37 CLK ICV_32 $T=-535 8960 1 270 $X=-1225 $Y=8080
X841 GND 4 199 38 CLK ICV_32 $T=-535 13600 1 270 $X=-1225 $Y=12720
X842 GND 3 200 32 CLK ICV_32 $T=-535 18240 1 270 $X=-1225 $Y=17360
X843 GND 2 201 33 CLK ICV_32 $T=-535 22880 1 270 $X=-1225 $Y=22000
X844 VDD 29 875 p18_CDNS_673871376604 $T=-9375 14680 0 270 $X=-9805 $Y=13945
X845 VDD A0 876 p18_CDNS_673871376604 $T=-9375 18300 0 270 $X=-9805 $Y=17565
X846 VDD 29 831 p18_CDNS_673871376604 $T=-9375 21920 0 270 $X=-9805 $Y=21185
X847 VDD A0 877 p18_CDNS_673871376604 $T=-9375 25540 0 270 $X=-9805 $Y=24805
X848 VDD 30 824 823 p18_CDNS_673871376603 $T=-9375 -230 0 270 $X=-9805 $Y=-965
X849 VDD A1 829 878 p18_CDNS_673871376603 $T=-9375 10630 0 270 $X=-9805 $Y=9895
X850 VDD 30 875 879 p18_CDNS_673871376603 $T=-9375 14250 0 270 $X=-9805 $Y=13515
X851 VDD 30 876 880 p18_CDNS_673871376603 $T=-9375 17870 0 270 $X=-9805 $Y=17135
X852 VDD A1 877 881 p18_CDNS_673871376603 $T=-9375 25110 0 270 $X=-9805 $Y=24375
X853 VDD 36 28 878 p18_CDNS_673871376602 $T=-9375 10200 0 270 $X=-9805 $Y=9110
X854 VDD 37 A2 879 p18_CDNS_673871376602 $T=-9375 13820 0 270 $X=-9805 $Y=12730
X855 VDD 38 A2 880 p18_CDNS_673871376602 $T=-9375 17440 0 270 $X=-9805 $Y=16350
X856 VDD 32 A2 830 p18_CDNS_673871376602 $T=-9375 21060 0 270 $X=-9805 $Y=19970
X857 VDD 33 A2 881 p18_CDNS_673871376602 $T=-9375 24680 0 270 $X=-9805 $Y=23590
X858 GND GND 28 A2 n18_CDNS_6738713766027 $T=-13045 -1400 1 270 $X=-13615 $Y=-2280
X859 GND GND 30 A1 n18_CDNS_6738713766027 $T=-13045 620 1 270 $X=-13615 $Y=-260
X860 GND 31 GND 28 n18_CDNS_6738713766027 $T=-11545 -1400 0 270 $X=-12685 $Y=-2280
X861 GND 34 GND A0 n18_CDNS_6738713766027 $T=-11545 3820 0 270 $X=-12685 $Y=2940
X862 GND 35 GND 28 n18_CDNS_6738713766027 $T=-11545 5840 0 270 $X=-12685 $Y=4960
X863 GND 35 GND 29 n18_CDNS_6738713766027 $T=-11545 7440 0 270 $X=-12685 $Y=6560
X864 GND 36 GND 28 n18_CDNS_6738713766027 $T=-11545 9460 0 270 $X=-12685 $Y=8580
X865 GND 36 GND A0 n18_CDNS_6738713766027 $T=-11545 11060 0 270 $X=-12685 $Y=10180
X866 GND 37 GND A2 n18_CDNS_6738713766027 $T=-11545 13080 0 270 $X=-12685 $Y=12200
X867 GND 37 GND 29 n18_CDNS_6738713766027 $T=-11545 14680 0 270 $X=-12685 $Y=13800
X868 GND 38 GND A2 n18_CDNS_6738713766027 $T=-11545 16700 0 270 $X=-12685 $Y=15820
X869 GND 38 GND A0 n18_CDNS_6738713766027 $T=-11545 18300 0 270 $X=-12685 $Y=17420
X870 GND 32 GND A2 n18_CDNS_6738713766027 $T=-11545 20320 0 270 $X=-12685 $Y=19440
X871 GND 32 GND 29 n18_CDNS_6738713766027 $T=-11545 21920 0 270 $X=-12685 $Y=21040
X872 GND 33 GND A2 n18_CDNS_6738713766027 $T=-11545 23940 0 270 $X=-12685 $Y=23060
X873 GND 33 GND A0 n18_CDNS_6738713766027 $T=-11545 25540 0 270 $X=-12685 $Y=24660
.ENDS
***************************************

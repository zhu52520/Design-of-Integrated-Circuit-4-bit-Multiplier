* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_672684331922 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672684331923 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 3 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672684331928 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=6 EP=5 IP=8 FDC=2
X0 1 2 4 6 p18_CDNS_672684331923 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 6 p18_CDNS_672684331928 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_672684331921 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672684331927 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672684331926 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6
** N=7 EP=6 IP=15 FDC=4
X0 1 5 7 n18_CDNS_672684331921 $T=0 0 0 0 $X=-660 $Y=-2020
X1 1 2 6 7 n18_CDNS_672684331927 $T=430 0 0 0 $X=110 $Y=-2020
X2 1 3 4 2 n18_CDNS_672684331926 $T=2370 0 0 0 $X=1710 $Y=-2020
X3 1 1 4 6 n18_CDNS_672684331926 $T=3810 0 0 0 $X=3150 $Y=-2020
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4
** N=4 EP=4 IP=8 FDC=2
X0 1 2 1 3 p18_CDNS_672684331922 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 1 4 p18_CDNS_672684331922 $T=1440 0 0 0 $X=530 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6726843319210 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X0 1 2 1 4 p18_CDNS_6726843319210 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 2 3 5 p18_CDNS_6726843319210 $T=1440 0 0 0 $X=530 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_6726843319211 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 3 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672684331929 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 3 6 n18_CDNS_672684331926 $T=-1950 0 0 0 $X=-2610 $Y=-2020
X1 1 4 5 6 n18_CDNS_672684331926 $T=0 0 0 0 $X=-660 $Y=-2020
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=3
X0 1 2 3 7 n18_CDNS_672684331926 $T=0 0 0 0 $X=-660 $Y=-2020
X1 1 4 5 6 7 8 ICV_5 $T=-2050 0 0 0 $X=-4660 $Y=-2020
.ENDS
***************************************
.SUBCKT n18_CDNS_672684331925 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 3 6 n18_CDNS_672684331925 $T=0 -1580 1 0 $X=-700 $Y=-2150
X1 1 4 5 6 n18_CDNS_672684331925 $T=0 0 0 0 $X=-700 $Y=-1180
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=4
X0 1 1 2 1 3 8 ICV_7 $T=0 0 0 0 $X=-700 $Y=-2150
X1 1 4 6 5 7 8 ICV_7 $T=2020 0 0 0 $X=1320 $Y=-2150
.ENDS
***************************************
.SUBCKT p18_CDNS_672684331920 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672684331924 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=4
X0 1 2 8 p18_CDNS_672684331920 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 8 p18_CDNS_672684331920 $T=0 2560 1 0 $X=-910 $Y=890
X2 1 4 5 2 p18_CDNS_672684331924 $T=2020 100 0 0 $X=1070 $Y=-430
X3 1 6 7 3 p18_CDNS_672684331924 $T=2020 2460 1 0 $X=1070 $Y=890
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=2
X0 1 2 5 p18_CDNS_672684331920 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 4 2 p18_CDNS_672684331924 $T=2020 100 0 0 $X=1070 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=4
X0 1 2 3 4 7 ICV_10 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 5 3 6 8 ICV_10 $T=4850 0 0 0 $X=3940 $Y=-430
.ENDS
***************************************
.SUBCKT vector_unit_v3 B3 X3 O8 O7 A3 A2 A1 A0 Y0 Y1 Y2 Y3 O6 O5 O4 O3 O2 O1 B2 X2
+ B1 X1 B0 X0 GND VDD O0
** N=489 EP=27 IP=1168 FDC=1178
M0 132 30 O8 GND NM L=1.8e-07 W=4.4e-07 $X=-20790 $Y=-27055 $D=0
M1 GND 141 6 GND NM L=1.8e-07 W=2.2e-07 $X=-20710 $Y=-52855 $D=0
M2 GND 10 3 GND NM L=1.8e-07 W=2.2e-07 $X=-20710 $Y=-49135 $D=0
M3 GND 11 4 GND NM L=1.8e-07 W=2.2e-07 $X=-20710 $Y=-1055 $D=0
M4 GND 142 7 GND NM L=1.8e-07 W=2.2e-07 $X=-20710 $Y=2665 $D=0
M5 GND 143 132 GND NM L=1.8e-07 W=4.4e-07 $X=-20070 $Y=-27055 $D=0
M6 10 15 19 GND NM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-40005 $D=0
M7 11 16 12 GND NM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-10405 $D=0
M8 GND 144 131 GND NM L=1.8e-07 W=4.4e-07 $X=-19870 $Y=-23355 $D=0
M9 143 19 GND GND NM L=1.8e-07 W=2.2e-07 $X=-19310 $Y=-26955 $D=0
M10 402 12 GND GND NM L=1.8e-07 W=4.4e-07 $X=-19150 $Y=-23355 $D=0
M11 144 19 402 GND NM L=1.8e-07 W=4.4e-07 $X=-18720 $Y=-23355 $D=0
M12 GND 133 17 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-68300 $D=0
M13 GND 134 8 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-66500 $D=0
M14 GND 135 59 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-61680 $D=0
M15 GND 136 77 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-59880 $D=0
M16 GND 137 79 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=9690 $D=0
M17 GND 138 60 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=11490 $D=0
M18 GND 139 9 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=16310 $D=0
M19 GND 140 18 GND NM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=18110 $D=0
M20 GND 8 156 GND NM L=1.8e-07 W=4.4e-07 $X=-16860 $Y=-52955 $D=0
M21 GND 6 157 GND NM L=1.8e-07 W=4.4e-07 $X=-16860 $Y=-49255 $D=0
M22 GND 7 158 GND NM L=1.8e-07 W=4.4e-07 $X=-16860 $Y=-1155 $D=0
M23 GND 9 159 GND NM L=1.8e-07 W=4.4e-07 $X=-16860 $Y=2545 $D=0
M24 173 144 155 GND NM L=1.8e-07 W=4.4e-07 $X=-16780 $Y=-23355 $D=0
M25 403 19 174 GND NM L=1.8e-07 W=4.4e-07 $X=-16530 $Y=-27055 $D=0
M26 163 48 15 GND NM L=1.8e-07 W=4.4e-07 $X=-16180 $Y=-36305 $D=0
M27 164 49 16 GND NM L=1.8e-07 W=4.4e-07 $X=-16180 $Y=-14105 $D=0
M28 GND 12 403 GND NM L=1.8e-07 W=4.4e-07 $X=-16100 $Y=-27055 $D=0
M29 GND 12 173 GND NM L=1.8e-07 W=4.4e-07 $X=-16060 $Y=-23355 $D=0
M30 GND 145 163 GND NM L=1.8e-07 W=4.4e-07 $X=-15460 $Y=-36305 $D=0
M31 GND 146 164 GND NM L=1.8e-07 W=4.4e-07 $X=-15460 $Y=-14105 $D=0
M32 174 143 GND GND NM L=1.8e-07 W=2.2e-07 $X=-15340 $Y=-26955 $D=0
M33 173 19 GND GND NM L=1.8e-07 W=4.4e-07 $X=-15340 $Y=-23355 $D=0
M34 GND 147 160 GND NM L=1.8e-07 W=4.4e-07 $X=-15260 $Y=-40005 $D=0
M35 GND 148 162 GND NM L=1.8e-07 W=4.4e-07 $X=-15260 $Y=-10405 $D=0
M36 145 24 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14700 $Y=-36185 $D=0
M37 146 25 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14700 $Y=-14005 $D=0
M38 404 20 GND GND NM L=1.8e-07 W=4.4e-07 $X=-14540 $Y=-40005 $D=0
M39 405 21 GND GND NM L=1.8e-07 W=4.4e-07 $X=-14540 $Y=-10405 $D=0
M40 33 149 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14160 $Y=-52855 $D=0
M41 20 150 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14160 $Y=-49135 $D=0
M42 21 151 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14160 $Y=-1055 $D=0
M43 34 152 GND GND NM L=1.8e-07 W=2.2e-07 $X=-14160 $Y=2665 $D=0
M44 147 24 404 GND NM L=1.8e-07 W=4.4e-07 $X=-14110 $Y=-40005 $D=0
M45 148 25 405 GND NM L=1.8e-07 W=4.4e-07 $X=-14110 $Y=-10405 $D=0
M46 175 174 GND GND NM L=1.8e-07 W=4.4e-07 $X=-13360 $Y=-27055 $D=0
M47 176 155 GND GND NM L=1.8e-07 W=4.4e-07 $X=-13360 $Y=-23355 $D=0
M48 GND 165 22 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-68300 $D=0
M49 GND 166 57 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-66500 $D=0
M50 GND 167 86 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-61680 $D=0
M51 GND 168 104 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-59880 $D=0
M52 GND 169 105 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=9690 $D=0
M53 GND 170 87 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=11490 $D=0
M54 GND 171 58 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=16310 $D=0
M55 GND 172 23 GND NM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=18110 $D=0
M56 O7 30 175 GND NM L=1.8e-07 W=4.4e-07 $X=-12600 $Y=-27055 $D=0
M57 GND 215 27 GND NM L=1.8e-07 W=4.4e-07 $X=-12180 $Y=-52955 $D=0
M58 GND 216 28 GND NM L=1.8e-07 W=4.4e-07 $X=-12180 $Y=2545 $D=0
M59 183 147 179 GND NM L=1.8e-07 W=4.4e-07 $X=-12170 $Y=-40005 $D=0
M60 184 148 180 GND NM L=1.8e-07 W=4.4e-07 $X=-12170 $Y=-10405 $D=0
M61 GND 185 24 GND NM L=1.8e-07 W=2.2e-07 $X=-12140 $Y=-49135 $D=0
M62 GND 186 25 GND NM L=1.8e-07 W=2.2e-07 $X=-12140 $Y=-1055 $D=0
M63 406 24 195 GND NM L=1.8e-07 W=4.4e-07 $X=-11920 $Y=-36305 $D=0
M64 407 25 196 GND NM L=1.8e-07 W=4.4e-07 $X=-11920 $Y=-14105 $D=0
M65 GND 20 406 GND NM L=1.8e-07 W=4.4e-07 $X=-11490 $Y=-36305 $D=0
M66 GND 21 407 GND NM L=1.8e-07 W=4.4e-07 $X=-11490 $Y=-14105 $D=0
M67 GND 20 183 GND NM L=1.8e-07 W=4.4e-07 $X=-11450 $Y=-40005 $D=0
M68 GND 21 184 GND NM L=1.8e-07 W=4.4e-07 $X=-11450 $Y=-10405 $D=0
M69 183 24 GND GND NM L=1.8e-07 W=4.4e-07 $X=-10730 $Y=-40005 $D=0
M70 195 145 GND GND NM L=1.8e-07 W=2.2e-07 $X=-10730 $Y=-36185 $D=0
M71 196 146 GND GND NM L=1.8e-07 W=2.2e-07 $X=-10730 $Y=-14005 $D=0
M72 184 25 GND GND NM L=1.8e-07 W=4.4e-07 $X=-10730 $Y=-10405 $D=0
M73 GND 59 208 GND NM L=1.8e-07 W=4.4e-07 $X=-10240 $Y=-52955 $D=0
M74 GND 60 209 GND NM L=1.8e-07 W=4.4e-07 $X=-10240 $Y=2545 $D=0
M75 408 59 GND GND NM L=1.8e-07 W=4.4e-07 $X=-9520 $Y=-52955 $D=0
M76 409 60 GND GND NM L=1.8e-07 W=4.4e-07 $X=-9520 $Y=2545 $D=0
M77 215 57 408 GND NM L=1.8e-07 W=4.4e-07 $X=-9090 $Y=-52955 $D=0
M78 216 58 409 GND NM L=1.8e-07 W=4.4e-07 $X=-9090 $Y=2545 $D=0
M79 201 179 GND GND NM L=1.8e-07 W=4.4e-07 $X=-8750 $Y=-40005 $D=0
M80 199 195 GND GND NM L=1.8e-07 W=4.4e-07 $X=-8750 $Y=-36305 $D=0
M81 200 196 GND GND NM L=1.8e-07 W=4.4e-07 $X=-8750 $Y=-14105 $D=0
M82 202 180 GND GND NM L=1.8e-07 W=4.4e-07 $X=-8750 $Y=-10405 $D=0
M83 204 65 30 GND NM L=1.8e-07 W=4.4e-07 $X=-8720 $Y=-27055 $D=0
M84 208 46 215 GND NM L=1.8e-07 W=4.4e-07 $X=-8370 $Y=-52955 $D=0
M85 209 47 216 GND NM L=1.8e-07 W=4.4e-07 $X=-8370 $Y=2545 $D=0
M86 GND 27 211 GND NM L=1.8e-07 W=4.4e-07 $X=-8290 $Y=-49255 $D=0
M87 GND 28 212 GND NM L=1.8e-07 W=4.4e-07 $X=-8290 $Y=-1155 $D=0
M88 GND 187 46 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-68300 $D=0
M89 GND 188 53 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-66500 $D=0
M90 GND 189 31 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-61680 $D=0
M91 GND 190 112 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-59880 $D=0
M92 GND 191 113 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=9690 $D=0
M93 GND 192 32 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=11490 $D=0
M94 GND 193 54 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=16310 $D=0
M95 GND 194 47 GND NM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=18110 $D=0
M96 GND 197 204 GND NM L=1.8e-07 W=4.4e-07 $X=-8000 $Y=-27055 $D=0
M97 52 48 199 GND NM L=1.8e-07 W=4.4e-07 $X=-7990 $Y=-36305 $D=0
M98 35 49 200 GND NM L=1.8e-07 W=4.4e-07 $X=-7990 $Y=-14105 $D=0
M99 GND 198 203 GND NM L=1.8e-07 W=4.4e-07 $X=-7800 $Y=-23355 $D=0
M100 GND 57 208 GND NM L=1.8e-07 W=4.4e-07 $X=-7650 $Y=-52955 $D=0
M101 GND 58 209 GND NM L=1.8e-07 W=4.4e-07 $X=-7650 $Y=2545 $D=0
M102 197 52 GND GND NM L=1.8e-07 W=2.2e-07 $X=-7240 $Y=-26955 $D=0
M103 410 35 GND GND NM L=1.8e-07 W=4.4e-07 $X=-7080 $Y=-23355 $D=0
M104 411 57 GND GND NM L=1.8e-07 W=4.4e-07 $X=-6930 $Y=-52955 $D=0
M105 412 58 GND GND NM L=1.8e-07 W=4.4e-07 $X=-6930 $Y=2545 $D=0
M106 198 52 410 GND NM L=1.8e-07 W=4.4e-07 $X=-6650 $Y=-23355 $D=0
M107 413 59 411 GND NM L=1.8e-07 W=4.4e-07 $X=-6500 $Y=-52955 $D=0
M108 414 60 412 GND NM L=1.8e-07 W=4.4e-07 $X=-6500 $Y=2545 $D=0
M109 240 46 413 GND NM L=1.8e-07 W=4.4e-07 $X=-6070 $Y=-52955 $D=0
M110 241 47 414 GND NM L=1.8e-07 W=4.4e-07 $X=-6070 $Y=2545 $D=0
M111 55 205 GND GND NM L=1.8e-07 W=2.2e-07 $X=-5590 $Y=-49135 $D=0
M112 56 206 GND GND NM L=1.8e-07 W=2.2e-07 $X=-5590 $Y=-1055 $D=0
M113 234 215 240 GND NM L=1.8e-07 W=4.4e-07 $X=-5350 $Y=-52955 $D=0
M114 235 216 241 GND NM L=1.8e-07 W=4.4e-07 $X=-5350 $Y=2545 $D=0
M115 239 198 229 GND NM L=1.8e-07 W=4.4e-07 $X=-4710 $Y=-23355 $D=0
M116 GND 46 234 GND NM L=1.8e-07 W=4.4e-07 $X=-4630 $Y=-52955 $D=0
M117 GND 47 235 GND NM L=1.8e-07 W=4.4e-07 $X=-4630 $Y=2545 $D=0
M118 415 52 242 GND NM L=1.8e-07 W=4.4e-07 $X=-4460 $Y=-27055 $D=0
M119 237 75 48 GND NM L=1.8e-07 W=4.4e-07 $X=-4110 $Y=-36305 $D=0
M120 238 76 49 GND NM L=1.8e-07 W=4.4e-07 $X=-4110 $Y=-14105 $D=0
M121 GND 35 415 GND NM L=1.8e-07 W=4.4e-07 $X=-4030 $Y=-27055 $D=0
M122 GND 35 239 GND NM L=1.8e-07 W=4.4e-07 $X=-3990 $Y=-23355 $D=0
M123 234 59 GND GND NM L=1.8e-07 W=4.4e-07 $X=-3910 $Y=-52955 $D=0
M124 235 60 GND GND NM L=1.8e-07 W=4.4e-07 $X=-3910 $Y=2545 $D=0
M125 GND 261 63 GND NM L=1.8e-07 W=4.4e-07 $X=-3610 $Y=-49255 $D=0
M126 GND 262 64 GND NM L=1.8e-07 W=4.4e-07 $X=-3610 $Y=-1155 $D=0
M127 GND 225 237 GND NM L=1.8e-07 W=4.4e-07 $X=-3390 $Y=-36305 $D=0
M128 GND 226 238 GND NM L=1.8e-07 W=4.4e-07 $X=-3390 $Y=-14105 $D=0
M129 GND 217 50 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-68300 $D=0
M130 GND 218 101 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-66500 $D=0
M131 GND 219 115 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-61680 $D=0
M132 GND 220 129 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-59880 $D=0
M133 GND 221 130 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=9690 $D=0
M134 GND 222 116 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=11490 $D=0
M135 GND 223 102 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=16310 $D=0
M136 GND 224 51 GND NM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=18110 $D=0
M137 242 197 GND GND NM L=1.8e-07 W=2.2e-07 $X=-3270 $Y=-26955 $D=0
M138 239 52 GND GND NM L=1.8e-07 W=4.4e-07 $X=-3270 $Y=-23355 $D=0
M139 GND 57 234 GND NM L=1.8e-07 W=4.4e-07 $X=-3190 $Y=-52955 $D=0
M140 GND 227 230 GND NM L=1.8e-07 W=4.4e-07 $X=-3190 $Y=-40005 $D=0
M141 GND 228 232 GND NM L=1.8e-07 W=4.4e-07 $X=-3190 $Y=-10405 $D=0
M142 GND 58 235 GND NM L=1.8e-07 W=4.4e-07 $X=-3190 $Y=2545 $D=0
M143 225 63 GND GND NM L=1.8e-07 W=2.2e-07 $X=-2630 $Y=-36185 $D=0
M144 226 64 GND GND NM L=1.8e-07 W=2.2e-07 $X=-2630 $Y=-14005 $D=0
M145 66 240 GND GND NM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=-52955 $D=0
M146 416 55 GND GND NM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=-40005 $D=0
M147 417 56 GND GND NM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=-10405 $D=0
M148 67 241 GND GND NM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=2545 $D=0
M149 227 63 416 GND NM L=1.8e-07 W=4.4e-07 $X=-2040 $Y=-40005 $D=0
M150 228 64 417 GND NM L=1.8e-07 W=4.4e-07 $X=-2040 $Y=-10405 $D=0
M151 GND 69 245 GND NM L=1.8e-07 W=4.4e-07 $X=-1670 $Y=-49255 $D=0
M152 GND 70 248 GND NM L=1.8e-07 W=4.4e-07 $X=-1670 $Y=-1155 $D=0
M153 243 242 GND GND NM L=1.8e-07 W=4.4e-07 $X=-1290 $Y=-27055 $D=0
M154 244 229 GND GND NM L=1.8e-07 W=4.4e-07 $X=-1290 $Y=-23355 $D=0
M155 418 69 GND GND NM L=1.8e-07 W=4.4e-07 $X=-950 $Y=-49255 $D=0
M156 419 70 GND GND NM L=1.8e-07 W=4.4e-07 $X=-950 $Y=-1155 $D=0
M157 O6 65 243 GND NM L=1.8e-07 W=4.4e-07 $X=-530 $Y=-27055 $D=0
M158 261 73 418 GND NM L=1.8e-07 W=4.4e-07 $X=-520 $Y=-49255 $D=0
M159 262 74 419 GND NM L=1.8e-07 W=4.4e-07 $X=-520 $Y=-1155 $D=0
M160 GND 253 73 GND NM L=1.8e-07 W=2.2e-07 $X=-490 $Y=-52855 $D=0
M161 GND 254 74 GND NM L=1.8e-07 W=2.2e-07 $X=-490 $Y=2665 $D=0
M162 255 227 249 GND NM L=1.8e-07 W=4.4e-07 $X=-100 $Y=-40005 $D=0
M163 256 228 250 GND NM L=1.8e-07 W=4.4e-07 $X=-100 $Y=-10405 $D=0
M164 420 63 257 GND NM L=1.8e-07 W=4.4e-07 $X=150 $Y=-36305 $D=0
M165 421 64 258 GND NM L=1.8e-07 W=4.4e-07 $X=150 $Y=-14105 $D=0
M166 245 66 261 GND NM L=1.8e-07 W=4.4e-07 $X=200 $Y=-49255 $D=0
M167 248 67 262 GND NM L=1.8e-07 W=4.4e-07 $X=200 $Y=-1155 $D=0
M168 GND 55 420 GND NM L=1.8e-07 W=4.4e-07 $X=580 $Y=-36305 $D=0
M169 GND 56 421 GND NM L=1.8e-07 W=4.4e-07 $X=580 $Y=-14105 $D=0
M170 GND 55 255 GND NM L=1.8e-07 W=4.4e-07 $X=620 $Y=-40005 $D=0
M171 GND 56 256 GND NM L=1.8e-07 W=4.4e-07 $X=620 $Y=-10405 $D=0
M172 GND 73 245 GND NM L=1.8e-07 W=4.4e-07 $X=920 $Y=-49255 $D=0
M173 GND 74 248 GND NM L=1.8e-07 W=4.4e-07 $X=920 $Y=-1155 $D=0
M174 255 63 GND GND NM L=1.8e-07 W=4.4e-07 $X=1340 $Y=-40005 $D=0
M175 257 225 GND GND NM L=1.8e-07 W=2.2e-07 $X=1340 $Y=-36185 $D=0
M176 258 226 GND GND NM L=1.8e-07 W=2.2e-07 $X=1340 $Y=-14005 $D=0
M177 256 64 GND GND NM L=1.8e-07 W=4.4e-07 $X=1340 $Y=-10405 $D=0
M178 422 73 GND GND NM L=1.8e-07 W=4.4e-07 $X=1640 $Y=-49255 $D=0
M179 423 74 GND GND NM L=1.8e-07 W=4.4e-07 $X=1640 $Y=-1155 $D=0
M180 424 69 422 GND NM L=1.8e-07 W=4.4e-07 $X=2070 $Y=-49255 $D=0
M181 425 70 423 GND NM L=1.8e-07 W=4.4e-07 $X=2070 $Y=-1155 $D=0
M182 277 66 424 GND NM L=1.8e-07 W=4.4e-07 $X=2500 $Y=-49255 $D=0
M183 278 67 425 GND NM L=1.8e-07 W=4.4e-07 $X=2500 $Y=-1155 $D=0
M184 273 261 277 GND NM L=1.8e-07 W=4.4e-07 $X=3220 $Y=-49255 $D=0
M185 276 262 278 GND NM L=1.8e-07 W=4.4e-07 $X=3220 $Y=-1155 $D=0
M186 267 249 GND GND NM L=1.8e-07 W=4.4e-07 $X=3320 $Y=-40005 $D=0
M187 265 257 GND GND NM L=1.8e-07 W=4.4e-07 $X=3320 $Y=-36305 $D=0
M188 266 258 GND GND NM L=1.8e-07 W=4.4e-07 $X=3320 $Y=-14105 $D=0
M189 268 250 GND GND NM L=1.8e-07 W=4.4e-07 $X=3320 $Y=-10405 $D=0
M190 270 88 65 GND NM L=1.8e-07 W=4.4e-07 $X=3350 $Y=-27055 $D=0
M191 GND 53 271 GND NM L=1.8e-07 W=4.4e-07 $X=3360 $Y=-52955 $D=0
M192 GND 54 272 GND NM L=1.8e-07 W=4.4e-07 $X=3360 $Y=2545 $D=0
M193 GND 66 273 GND NM L=1.8e-07 W=4.4e-07 $X=3940 $Y=-49255 $D=0
M194 GND 67 276 GND NM L=1.8e-07 W=4.4e-07 $X=3940 $Y=-1155 $D=0
M195 GND 259 270 GND NM L=1.8e-07 W=4.4e-07 $X=4070 $Y=-27055 $D=0
M196 78 75 265 GND NM L=1.8e-07 W=4.4e-07 $X=4080 $Y=-36305 $D=0
M197 68 76 266 GND NM L=1.8e-07 W=4.4e-07 $X=4080 $Y=-14105 $D=0
M198 GND 260 269 GND NM L=1.8e-07 W=4.4e-07 $X=4270 $Y=-23355 $D=0
M199 273 69 GND GND NM L=1.8e-07 W=4.4e-07 $X=4660 $Y=-49255 $D=0
M200 276 70 GND GND NM L=1.8e-07 W=4.4e-07 $X=4660 $Y=-1155 $D=0
M201 259 78 GND GND NM L=1.8e-07 W=2.2e-07 $X=4830 $Y=-26955 $D=0
M202 426 68 GND GND NM L=1.8e-07 W=4.4e-07 $X=4990 $Y=-23355 $D=0
M203 GND 73 273 GND NM L=1.8e-07 W=4.4e-07 $X=5380 $Y=-49255 $D=0
M204 GND 74 276 GND NM L=1.8e-07 W=4.4e-07 $X=5380 $Y=-1155 $D=0
M205 260 78 426 GND NM L=1.8e-07 W=4.4e-07 $X=5420 $Y=-23355 $D=0
M206 93 263 GND GND NM L=1.8e-07 W=2.2e-07 $X=6060 $Y=-52855 $D=0
M207 94 264 GND GND NM L=1.8e-07 W=2.2e-07 $X=6060 $Y=2665 $D=0
M208 80 277 GND GND NM L=1.8e-07 W=4.4e-07 $X=6100 $Y=-49255 $D=0
M209 81 278 GND GND NM L=1.8e-07 W=4.4e-07 $X=6100 $Y=-1155 $D=0
M210 293 260 287 GND NM L=1.8e-07 W=4.4e-07 $X=7360 $Y=-23355 $D=0
M211 427 78 294 GND NM L=1.8e-07 W=4.4e-07 $X=7610 $Y=-27055 $D=0
M212 291 285 75 GND NM L=1.8e-07 W=4.4e-07 $X=7960 $Y=-36305 $D=0
M213 292 286 76 GND NM L=1.8e-07 W=4.4e-07 $X=7960 $Y=-14105 $D=0
M214 GND 317 82 GND NM L=1.8e-07 W=4.4e-07 $X=8040 $Y=-49255 $D=0
M215 GND 68 427 GND NM L=1.8e-07 W=4.4e-07 $X=8040 $Y=-27055 $D=0
M216 GND 318 83 GND NM L=1.8e-07 W=4.4e-07 $X=8040 $Y=-1155 $D=0
M217 GND 295 69 GND NM L=1.8e-07 W=2.2e-07 $X=8080 $Y=-52855 $D=0
M218 GND 68 293 GND NM L=1.8e-07 W=4.4e-07 $X=8080 $Y=-23355 $D=0
M219 GND 296 70 GND NM L=1.8e-07 W=2.2e-07 $X=8080 $Y=2665 $D=0
M220 GND 279 291 GND NM L=1.8e-07 W=4.4e-07 $X=8680 $Y=-36305 $D=0
M221 GND 280 292 GND NM L=1.8e-07 W=4.4e-07 $X=8680 $Y=-14105 $D=0
M222 294 259 GND GND NM L=1.8e-07 W=2.2e-07 $X=8800 $Y=-26955 $D=0
M223 293 78 GND GND NM L=1.8e-07 W=4.4e-07 $X=8800 $Y=-23355 $D=0
M224 GND 281 288 GND NM L=1.8e-07 W=4.4e-07 $X=8880 $Y=-40005 $D=0
M225 GND 282 290 GND NM L=1.8e-07 W=4.4e-07 $X=8880 $Y=-10405 $D=0
M226 279 82 GND GND NM L=1.8e-07 W=2.2e-07 $X=9440 $Y=-36185 $D=0
M227 280 83 GND GND NM L=1.8e-07 W=2.2e-07 $X=9440 $Y=-14005 $D=0
M228 428 80 GND GND NM L=1.8e-07 W=4.4e-07 $X=9600 $Y=-40005 $D=0
M229 429 81 GND GND NM L=1.8e-07 W=4.4e-07 $X=9600 $Y=-10405 $D=0
M230 GND 91 301 GND NM L=1.8e-07 W=4.4e-07 $X=9980 $Y=-49255 $D=0
M231 GND 92 304 GND NM L=1.8e-07 W=4.4e-07 $X=9980 $Y=-1155 $D=0
M232 281 82 428 GND NM L=1.8e-07 W=4.4e-07 $X=10030 $Y=-40005 $D=0
M233 282 83 429 GND NM L=1.8e-07 W=4.4e-07 $X=10030 $Y=-10405 $D=0
M234 430 91 GND GND NM L=1.8e-07 W=4.4e-07 $X=10700 $Y=-49255 $D=0
M235 431 92 GND GND NM L=1.8e-07 W=4.4e-07 $X=10700 $Y=-1155 $D=0
M236 297 294 GND GND NM L=1.8e-07 W=4.4e-07 $X=10780 $Y=-27055 $D=0
M237 298 287 GND GND NM L=1.8e-07 W=4.4e-07 $X=10780 $Y=-23355 $D=0
M238 317 93 430 GND NM L=1.8e-07 W=4.4e-07 $X=11130 $Y=-49255 $D=0
M239 318 94 431 GND NM L=1.8e-07 W=4.4e-07 $X=11130 $Y=-1155 $D=0
M240 O5 88 297 GND NM L=1.8e-07 W=4.4e-07 $X=11540 $Y=-27055 $D=0
M241 301 89 317 GND NM L=1.8e-07 W=4.4e-07 $X=11850 $Y=-49255 $D=0
M242 304 90 318 GND NM L=1.8e-07 W=4.4e-07 $X=11850 $Y=-1155 $D=0
M243 GND 77 307 GND NM L=1.8e-07 W=4.4e-07 $X=11930 $Y=-52955 $D=0
M244 GND 79 308 GND NM L=1.8e-07 W=4.4e-07 $X=11930 $Y=2545 $D=0
M245 311 281 305 GND NM L=1.8e-07 W=4.4e-07 $X=11970 $Y=-40005 $D=0
M246 312 282 306 GND NM L=1.8e-07 W=4.4e-07 $X=11970 $Y=-10405 $D=0
M247 432 82 313 GND NM L=1.8e-07 W=4.4e-07 $X=12220 $Y=-36305 $D=0
M248 433 83 314 GND NM L=1.8e-07 W=4.4e-07 $X=12220 $Y=-14105 $D=0
M249 GND 93 301 GND NM L=1.8e-07 W=4.4e-07 $X=12570 $Y=-49255 $D=0
M250 GND 94 304 GND NM L=1.8e-07 W=4.4e-07 $X=12570 $Y=-1155 $D=0
M251 GND 80 432 GND NM L=1.8e-07 W=4.4e-07 $X=12650 $Y=-36305 $D=0
M252 GND 81 433 GND NM L=1.8e-07 W=4.4e-07 $X=12650 $Y=-14105 $D=0
M253 GND 80 311 GND NM L=1.8e-07 W=4.4e-07 $X=12690 $Y=-40005 $D=0
M254 GND 81 312 GND NM L=1.8e-07 W=4.4e-07 $X=12690 $Y=-10405 $D=0
M255 434 93 GND GND NM L=1.8e-07 W=4.4e-07 $X=13290 $Y=-49255 $D=0
M256 435 94 GND GND NM L=1.8e-07 W=4.4e-07 $X=13290 $Y=-1155 $D=0
M257 311 82 GND GND NM L=1.8e-07 W=4.4e-07 $X=13410 $Y=-40005 $D=0
M258 313 279 GND GND NM L=1.8e-07 W=2.2e-07 $X=13410 $Y=-36185 $D=0
M259 314 280 GND GND NM L=1.8e-07 W=2.2e-07 $X=13410 $Y=-14005 $D=0
M260 312 83 GND GND NM L=1.8e-07 W=4.4e-07 $X=13410 $Y=-10405 $D=0
M261 436 91 434 GND NM L=1.8e-07 W=4.4e-07 $X=13720 $Y=-49255 $D=0
M262 437 92 435 GND NM L=1.8e-07 W=4.4e-07 $X=13720 $Y=-1155 $D=0
M263 329 89 436 GND NM L=1.8e-07 W=4.4e-07 $X=14150 $Y=-49255 $D=0
M264 330 90 437 GND NM L=1.8e-07 W=4.4e-07 $X=14150 $Y=-1155 $D=0
M265 91 299 GND GND NM L=1.8e-07 W=2.2e-07 $X=14630 $Y=-52855 $D=0
M266 92 300 GND GND NM L=1.8e-07 W=2.2e-07 $X=14630 $Y=2665 $D=0
M267 325 317 329 GND NM L=1.8e-07 W=4.4e-07 $X=14870 $Y=-49255 $D=0
M268 328 318 330 GND NM L=1.8e-07 W=4.4e-07 $X=14870 $Y=-1155 $D=0
M269 321 305 GND GND NM L=1.8e-07 W=4.4e-07 $X=15390 $Y=-40005 $D=0
M270 319 313 GND GND NM L=1.8e-07 W=4.4e-07 $X=15390 $Y=-36305 $D=0
M271 320 314 GND GND NM L=1.8e-07 W=4.4e-07 $X=15390 $Y=-14105 $D=0
M272 322 306 GND GND NM L=1.8e-07 W=4.4e-07 $X=15390 $Y=-10405 $D=0
M273 324 109 88 GND NM L=1.8e-07 W=4.4e-07 $X=15420 $Y=-27055 $D=0
M274 GND 89 325 GND NM L=1.8e-07 W=4.4e-07 $X=15590 $Y=-49255 $D=0
M275 GND 90 328 GND NM L=1.8e-07 W=4.4e-07 $X=15590 $Y=-1155 $D=0
M276 GND 315 324 GND NM L=1.8e-07 W=4.4e-07 $X=16140 $Y=-27055 $D=0
M277 98 285 319 GND NM L=1.8e-07 W=4.4e-07 $X=16150 $Y=-36305 $D=0
M278 95 286 320 GND NM L=1.8e-07 W=4.4e-07 $X=16150 $Y=-14105 $D=0
M279 325 91 GND GND NM L=1.8e-07 W=4.4e-07 $X=16310 $Y=-49255 $D=0
M280 328 92 GND GND NM L=1.8e-07 W=4.4e-07 $X=16310 $Y=-1155 $D=0
M281 GND 316 323 GND NM L=1.8e-07 W=4.4e-07 $X=16340 $Y=-23355 $D=0
M282 GND 347 89 GND NM L=1.8e-07 W=4.4e-07 $X=16610 $Y=-52955 $D=0
M283 GND 348 90 GND NM L=1.8e-07 W=4.4e-07 $X=16610 $Y=2545 $D=0
M284 315 98 GND GND NM L=1.8e-07 W=2.2e-07 $X=16900 $Y=-26955 $D=0
M285 GND 93 325 GND NM L=1.8e-07 W=4.4e-07 $X=17030 $Y=-49255 $D=0
M286 GND 94 328 GND NM L=1.8e-07 W=4.4e-07 $X=17030 $Y=-1155 $D=0
M287 438 95 GND GND NM L=1.8e-07 W=4.4e-07 $X=17060 $Y=-23355 $D=0
M288 316 98 438 GND NM L=1.8e-07 W=4.4e-07 $X=17490 $Y=-23355 $D=0
M289 99 329 GND GND NM L=1.8e-07 W=4.4e-07 $X=17750 $Y=-49255 $D=0
M290 100 330 GND GND NM L=1.8e-07 W=4.4e-07 $X=17750 $Y=-1155 $D=0
M291 GND 283 285 GND NM L=1.8e-07 W=2.2e-07 $X=18130 $Y=-39905 $D=0
M292 GND 284 286 GND NM L=1.8e-07 W=2.2e-07 $X=18130 $Y=-10285 $D=0
M293 GND 104 334 GND NM L=1.8e-07 W=4.4e-07 $X=18550 $Y=-52955 $D=0
M294 GND 105 335 GND NM L=1.8e-07 W=4.4e-07 $X=18550 $Y=2545 $D=0
M295 439 104 GND GND NM L=1.8e-07 W=4.4e-07 $X=19270 $Y=-52955 $D=0
M296 440 105 GND GND NM L=1.8e-07 W=4.4e-07 $X=19270 $Y=2545 $D=0
M297 337 316 331 GND NM L=1.8e-07 W=4.4e-07 $X=19430 $Y=-23355 $D=0
M298 441 98 338 GND NM L=1.8e-07 W=4.4e-07 $X=19680 $Y=-27055 $D=0
M299 347 31 439 GND NM L=1.8e-07 W=4.4e-07 $X=19700 $Y=-52955 $D=0
M300 348 32 440 GND NM L=1.8e-07 W=4.4e-07 $X=19700 $Y=2545 $D=0
M301 GND 339 96 GND NM L=1.8e-07 W=2.2e-07 $X=19730 $Y=-49135 $D=0
M302 GND 340 97 GND NM L=1.8e-07 W=2.2e-07 $X=19730 $Y=-1055 $D=0
M303 GND 95 441 GND NM L=1.8e-07 W=4.4e-07 $X=20110 $Y=-27055 $D=0
M304 GND 95 337 GND NM L=1.8e-07 W=4.4e-07 $X=20150 $Y=-23355 $D=0
M305 334 101 347 GND NM L=1.8e-07 W=4.4e-07 $X=20420 $Y=-52955 $D=0
M306 335 102 348 GND NM L=1.8e-07 W=4.4e-07 $X=20420 $Y=2545 $D=0
M307 338 315 GND GND NM L=1.8e-07 W=2.2e-07 $X=20870 $Y=-26955 $D=0
M308 337 98 GND GND NM L=1.8e-07 W=4.4e-07 $X=20870 $Y=-23355 $D=0
M309 GND 31 334 GND NM L=1.8e-07 W=4.4e-07 $X=21140 $Y=-52955 $D=0
M310 GND 32 335 GND NM L=1.8e-07 W=4.4e-07 $X=21140 $Y=2545 $D=0
M311 442 31 GND GND NM L=1.8e-07 W=4.4e-07 $X=21860 $Y=-52955 $D=0
M312 443 32 GND GND NM L=1.8e-07 W=4.4e-07 $X=21860 $Y=2545 $D=0
M313 GND 96 343 GND NM L=1.8e-07 W=4.4e-07 $X=21980 $Y=-40005 $D=0
M314 GND 97 344 GND NM L=1.8e-07 W=4.4e-07 $X=21980 $Y=-10405 $D=0
M315 444 104 442 GND NM L=1.8e-07 W=4.4e-07 $X=22290 $Y=-52955 $D=0
M316 445 105 443 GND NM L=1.8e-07 W=4.4e-07 $X=22290 $Y=2545 $D=0
M317 357 101 444 GND NM L=1.8e-07 W=4.4e-07 $X=22720 $Y=-52955 $D=0
M318 358 102 445 GND NM L=1.8e-07 W=4.4e-07 $X=22720 $Y=2545 $D=0
M319 345 338 GND GND NM L=1.8e-07 W=4.4e-07 $X=22850 $Y=-27055 $D=0
M320 346 331 GND GND NM L=1.8e-07 W=4.4e-07 $X=22850 $Y=-23355 $D=0
M321 354 347 357 GND NM L=1.8e-07 W=4.4e-07 $X=23440 $Y=-52955 $D=0
M322 355 348 358 GND NM L=1.8e-07 W=4.4e-07 $X=23440 $Y=2545 $D=0
M323 GND 110 351 GND NM L=1.8e-07 W=4.4e-07 $X=23580 $Y=-49255 $D=0
M324 GND 111 352 GND NM L=1.8e-07 W=4.4e-07 $X=23580 $Y=-1155 $D=0
M325 O4 109 345 GND NM L=1.8e-07 W=4.4e-07 $X=23610 $Y=-27055 $D=0
M326 GND 101 354 GND NM L=1.8e-07 W=4.4e-07 $X=24160 $Y=-52955 $D=0
M327 GND 102 355 GND NM L=1.8e-07 W=4.4e-07 $X=24160 $Y=2545 $D=0
M328 117 341 GND GND NM L=1.8e-07 W=2.2e-07 $X=24680 $Y=-39905 $D=0
M329 114 342 GND GND NM L=1.8e-07 W=2.2e-07 $X=24680 $Y=-10285 $D=0
M330 354 104 GND GND NM L=1.8e-07 W=4.4e-07 $X=24880 $Y=-52955 $D=0
M331 355 105 GND GND NM L=1.8e-07 W=4.4e-07 $X=24880 $Y=2545 $D=0
M332 GND 31 354 GND NM L=1.8e-07 W=4.4e-07 $X=25600 $Y=-52955 $D=0
M333 GND 32 355 GND NM L=1.8e-07 W=4.4e-07 $X=25600 $Y=2545 $D=0
M334 122 349 GND GND NM L=1.8e-07 W=2.2e-07 $X=26280 $Y=-49135 $D=0
M335 121 350 GND GND NM L=1.8e-07 W=2.2e-07 $X=26280 $Y=-1055 $D=0
M336 107 357 GND GND NM L=1.8e-07 W=4.4e-07 $X=26320 $Y=-52955 $D=0
M337 108 358 GND GND NM L=1.8e-07 W=4.4e-07 $X=26320 $Y=2545 $D=0
M338 362 120 109 GND NM L=1.8e-07 W=4.4e-07 $X=27490 $Y=-27055 $D=0
M339 GND 359 362 GND NM L=1.8e-07 W=4.4e-07 $X=28210 $Y=-27055 $D=0
M340 GND 363 110 GND NM L=1.8e-07 W=2.2e-07 $X=28300 $Y=-52855 $D=0
M341 GND 364 111 GND NM L=1.8e-07 W=2.2e-07 $X=28300 $Y=2665 $D=0
M342 GND 360 361 GND NM L=1.8e-07 W=4.4e-07 $X=28410 $Y=-23355 $D=0
M343 359 117 GND GND NM L=1.8e-07 W=2.2e-07 $X=28970 $Y=-26955 $D=0
M344 446 114 GND GND NM L=1.8e-07 W=4.4e-07 $X=29130 $Y=-23355 $D=0
M345 360 117 446 GND NM L=1.8e-07 W=4.4e-07 $X=29560 $Y=-23355 $D=0
M346 371 360 367 GND NM L=1.8e-07 W=4.4e-07 $X=31500 $Y=-23355 $D=0
M347 447 117 372 GND NM L=1.8e-07 W=4.4e-07 $X=31750 $Y=-27055 $D=0
M348 GND 112 369 GND NM L=1.8e-07 W=4.4e-07 $X=32150 $Y=-52955 $D=0
M349 GND 113 370 GND NM L=1.8e-07 W=4.4e-07 $X=32150 $Y=2545 $D=0
M350 GND 114 447 GND NM L=1.8e-07 W=4.4e-07 $X=32180 $Y=-27055 $D=0
M351 GND 114 371 GND NM L=1.8e-07 W=4.4e-07 $X=32220 $Y=-23355 $D=0
M352 372 359 GND GND NM L=1.8e-07 W=2.2e-07 $X=32940 $Y=-26955 $D=0
M353 371 117 GND GND NM L=1.8e-07 W=4.4e-07 $X=32940 $Y=-23355 $D=0
M354 127 365 GND GND NM L=1.8e-07 W=2.2e-07 $X=34850 $Y=-52855 $D=0
M355 126 366 GND GND NM L=1.8e-07 W=2.2e-07 $X=34850 $Y=2665 $D=0
M356 373 372 GND GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=-27055 $D=0
M357 374 367 GND GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=-23355 $D=0
M358 O3 120 373 GND NM L=1.8e-07 W=4.4e-07 $X=35680 $Y=-27055 $D=0
M359 378 125 120 GND NM L=1.8e-07 W=4.4e-07 $X=39560 $Y=-27055 $D=0
M360 GND 375 378 GND NM L=1.8e-07 W=4.4e-07 $X=40280 $Y=-27055 $D=0
M361 GND 376 377 GND NM L=1.8e-07 W=4.4e-07 $X=40480 $Y=-23355 $D=0
M362 375 122 GND GND NM L=1.8e-07 W=2.2e-07 $X=41040 $Y=-26955 $D=0
M363 448 121 GND GND NM L=1.8e-07 W=4.4e-07 $X=41200 $Y=-23355 $D=0
M364 376 122 448 GND NM L=1.8e-07 W=4.4e-07 $X=41630 $Y=-23355 $D=0
M365 381 376 379 GND NM L=1.8e-07 W=4.4e-07 $X=43570 $Y=-23355 $D=0
M366 449 122 382 GND NM L=1.8e-07 W=4.4e-07 $X=43820 $Y=-27055 $D=0
M367 GND 121 449 GND NM L=1.8e-07 W=4.4e-07 $X=44250 $Y=-27055 $D=0
M368 GND 121 381 GND NM L=1.8e-07 W=4.4e-07 $X=44290 $Y=-23355 $D=0
M369 382 375 GND GND NM L=1.8e-07 W=2.2e-07 $X=45010 $Y=-26955 $D=0
M370 381 122 GND GND NM L=1.8e-07 W=4.4e-07 $X=45010 $Y=-23355 $D=0
M371 383 382 GND GND NM L=1.8e-07 W=4.4e-07 $X=46990 $Y=-27055 $D=0
M372 384 379 GND GND NM L=1.8e-07 W=4.4e-07 $X=46990 $Y=-23355 $D=0
M373 O2 125 383 GND NM L=1.8e-07 W=4.4e-07 $X=47750 $Y=-27055 $D=0
M374 390 388 125 GND NM L=1.8e-07 W=4.4e-07 $X=51630 $Y=-27055 $D=0
M375 GND 385 390 GND NM L=1.8e-07 W=4.4e-07 $X=52350 $Y=-27055 $D=0
M376 GND 386 389 GND NM L=1.8e-07 W=4.4e-07 $X=52550 $Y=-23355 $D=0
M377 385 127 GND GND NM L=1.8e-07 W=2.2e-07 $X=53110 $Y=-26955 $D=0
M378 450 126 GND GND NM L=1.8e-07 W=4.4e-07 $X=53270 $Y=-23355 $D=0
M379 386 127 450 GND NM L=1.8e-07 W=4.4e-07 $X=53700 $Y=-23355 $D=0
M380 393 386 391 GND NM L=1.8e-07 W=4.4e-07 $X=55640 $Y=-23355 $D=0
M381 451 127 394 GND NM L=1.8e-07 W=4.4e-07 $X=55890 $Y=-27055 $D=0
M382 GND 126 451 GND NM L=1.8e-07 W=4.4e-07 $X=56320 $Y=-27055 $D=0
M383 GND 126 393 GND NM L=1.8e-07 W=4.4e-07 $X=56360 $Y=-23355 $D=0
M384 394 385 GND GND NM L=1.8e-07 W=2.2e-07 $X=57080 $Y=-26955 $D=0
M385 393 127 GND GND NM L=1.8e-07 W=4.4e-07 $X=57080 $Y=-23355 $D=0
M386 395 394 GND GND NM L=1.8e-07 W=4.4e-07 $X=59060 $Y=-27055 $D=0
M387 396 391 GND GND NM L=1.8e-07 W=4.4e-07 $X=59060 $Y=-23355 $D=0
M388 O1 388 395 GND NM L=1.8e-07 W=4.4e-07 $X=59820 $Y=-27055 $D=0
M389 GND 387 388 GND NM L=1.8e-07 W=2.2e-07 $X=61800 $Y=-23235 $D=0
M390 GND 129 398 GND NM L=1.8e-07 W=4.4e-07 $X=65650 $Y=-23355 $D=0
M391 O0 397 GND GND NM L=1.8e-07 W=2.2e-07 $X=68350 $Y=-23235 $D=0
M392 131 30 O8 VDD PM L=1.8e-07 W=4.4e-07 $X=-20670 $Y=-19910 $D=4
M393 141 8 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-56400 $D=4
M394 10 6 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-45810 $D=4
M395 10 13 19 VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-43450 $D=4
M396 11 14 12 VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-6960 $D=4
M397 11 7 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=-4600 $D=4
M398 142 9 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-19950 $Y=5990 $D=4
M399 VDD 143 132 VDD PM L=1.8e-07 W=8.8e-07 $X=-19870 $Y=-30500 $D=4
M400 144 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-19150 $Y=-19910 $D=4
M401 143 12 452 VDD PM L=1.8e-07 W=8.8e-07 $X=-18720 $Y=-30500 $D=4
M402 77 136 A0 VDD PM L=1.8e-07 W=2.2e-07 $X=-18650 $Y=-58540 $D=4
M403 79 137 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=-18650 $Y=8350 $D=4
M404 VDD 19 144 VDD PM L=1.8e-07 W=4.4e-07 $X=-18430 $Y=-19910 $D=4
M405 GND B3 17 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-69640 $D=4
M406 GND B3 8 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-65160 $D=4
M407 GND B3 59 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-63020 $D=4
M408 GND B3 77 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=-58540 $D=4
M409 GND X3 79 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=8350 $D=4
M410 GND X3 60 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=12830 $D=4
M411 GND X3 9 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=14970 $D=4
M412 GND X3 18 VDD PM L=1.8e-07 W=2.2e-07 $X=-17850 $Y=19450 $D=4
M413 149 141 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-17290 $Y=-56400 $D=4
M414 150 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-17290 $Y=-45810 $D=4
M415 151 11 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-17290 $Y=-4600 $D=4
M416 152 142 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-17290 $Y=5990 $D=4
M417 155 144 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-16490 $Y=-19910 $D=4
M418 VDD 17 453 VDD PM L=1.8e-07 W=8.8e-07 $X=-16100 $Y=-46250 $D=4
M419 VDD 18 454 VDD PM L=1.8e-07 W=8.8e-07 $X=-16100 $Y=-4600 $D=4
M420 160 48 15 VDD PM L=1.8e-07 W=4.4e-07 $X=-16060 $Y=-43450 $D=4
M421 161 12 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-16060 $Y=-30500 $D=4
M422 162 49 16 VDD PM L=1.8e-07 W=4.4e-07 $X=-16060 $Y=-6960 $D=4
M423 163 36 15 VDD PM L=1.8e-07 W=4.4e-07 $X=-16020 $Y=-32860 $D=4
M424 168 B2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-15820 $Y=-58640 $D=4
M425 169 X2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-15820 $Y=8230 $D=4
M426 455 12 155 VDD PM L=1.8e-07 W=8.8e-07 $X=-15730 $Y=-20350 $D=4
M427 174 143 161 VDD PM L=1.8e-07 W=8.8e-07 $X=-15340 $Y=-30500 $D=4
M428 VDD 145 163 VDD PM L=1.8e-07 W=8.8e-07 $X=-15260 $Y=-33300 $D=4
M429 VDD 146 164 VDD PM L=1.8e-07 W=8.8e-07 $X=-15260 $Y=-17550 $D=4
M430 147 20 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-14540 $Y=-43450 $D=4
M431 456 25 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-14540 $Y=-17550 $D=4
M432 148 21 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-14540 $Y=-6960 $D=4
M433 145 20 457 VDD PM L=1.8e-07 W=8.8e-07 $X=-14110 $Y=-33300 $D=4
M434 VDD 24 147 VDD PM L=1.8e-07 W=4.4e-07 $X=-13820 $Y=-43450 $D=4
M435 VDD 25 148 VDD PM L=1.8e-07 W=4.4e-07 $X=-13820 $Y=-6960 $D=4
M436 104 168 A0 VDD PM L=1.8e-07 W=2.2e-07 $X=-13800 $Y=-58540 $D=4
M437 105 169 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=-13800 $Y=8350 $D=4
M438 176 155 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-13360 $Y=-20350 $D=4
M439 GND B2 22 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-69640 $D=4
M440 GND B2 57 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-65160 $D=4
M441 GND B2 86 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-63020 $D=4
M442 GND B2 104 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=-58540 $D=4
M443 GND X2 105 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=8350 $D=4
M444 GND X2 87 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=12830 $D=4
M445 GND X2 58 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=14970 $D=4
M446 GND X2 23 VDD PM L=1.8e-07 W=2.2e-07 $X=-13000 $Y=19450 $D=4
M447 O7 29 175 VDD PM L=1.8e-07 W=4.4e-07 $X=-12640 $Y=-30500 $D=4
M448 O7 30 176 VDD PM L=1.8e-07 W=4.4e-07 $X=-12600 $Y=-19910 $D=4
M449 VDD 215 27 VDD PM L=1.8e-07 W=8.8e-07 $X=-12180 $Y=-56400 $D=4
M450 VDD 216 28 VDD PM L=1.8e-07 W=8.8e-07 $X=-12180 $Y=5550 $D=4
M451 VDD 24 181 VDD PM L=1.8e-07 W=8.8e-07 $X=-12170 $Y=-33300 $D=4
M452 179 147 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-11880 $Y=-43450 $D=4
M453 180 148 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-11880 $Y=-6960 $D=4
M454 181 20 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-11450 $Y=-33300 $D=4
M455 182 21 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-11450 $Y=-17550 $D=4
M456 185 27 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-11380 $Y=-45810 $D=4
M457 186 28 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-11380 $Y=-4600 $D=4
M458 VDD 24 458 VDD PM L=1.8e-07 W=8.8e-07 $X=-10690 $Y=-43450 $D=4
M459 VDD 25 459 VDD PM L=1.8e-07 W=8.8e-07 $X=-10690 $Y=-7400 $D=4
M460 VDD 33 185 VDD PM L=1.8e-07 W=4.4e-07 $X=-10660 $Y=-45810 $D=4
M461 VDD 34 186 VDD PM L=1.8e-07 W=4.4e-07 $X=-10660 $Y=-4600 $D=4
M462 198 65 29 VDD PM L=1.8e-07 W=4.4e-07 $X=-10550 $Y=-19910 $D=4
M463 197 62 29 VDD PM L=1.8e-07 W=4.4e-07 $X=-10500 $Y=-30500 $D=4
M464 VDD 59 207 VDD PM L=1.8e-07 W=8.8e-07 $X=-10240 $Y=-56400 $D=4
M465 VDD 60 210 VDD PM L=1.8e-07 W=8.8e-07 $X=-10240 $Y=5550 $D=4
M466 460 59 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-9520 $Y=-56400 $D=4
M467 461 60 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-9520 $Y=5550 $D=4
M468 215 57 460 VDD PM L=1.8e-07 W=8.8e-07 $X=-9090 $Y=-56400 $D=4
M469 216 58 461 VDD PM L=1.8e-07 W=8.8e-07 $X=-9090 $Y=5550 $D=4
M470 199 195 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-8790 $Y=-33300 $D=4
M471 200 196 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-8790 $Y=-17550 $D=4
M472 201 179 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-8750 $Y=-43450 $D=4
M473 202 180 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-8750 $Y=-7400 $D=4
M474 205 185 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-8720 $Y=-45810 $D=4
M475 206 186 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-8720 $Y=-4600 $D=4
M476 203 65 30 VDD PM L=1.8e-07 W=4.4e-07 $X=-8600 $Y=-19910 $D=4
M477 207 46 215 VDD PM L=1.8e-07 W=8.8e-07 $X=-8370 $Y=-56400 $D=4
M478 210 47 216 VDD PM L=1.8e-07 W=8.8e-07 $X=-8370 $Y=5550 $D=4
M479 GND B1 46 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-69640 $D=4
M480 GND B1 53 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-65160 $D=4
M481 GND B1 31 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-63020 $D=4
M482 GND B1 112 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=-58540 $D=4
M483 GND X1 113 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=8350 $D=4
M484 GND X1 32 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=12830 $D=4
M485 GND X1 54 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=14970 $D=4
M486 GND X1 47 VDD PM L=1.8e-07 W=2.2e-07 $X=-8150 $Y=19450 $D=4
M487 52 36 199 VDD PM L=1.8e-07 W=4.4e-07 $X=-8030 $Y=-32860 $D=4
M488 35 37 200 VDD PM L=1.8e-07 W=4.4e-07 $X=-8030 $Y=-17550 $D=4
M489 52 48 201 VDD PM L=1.8e-07 W=4.4e-07 $X=-7990 $Y=-43450 $D=4
M490 35 49 202 VDD PM L=1.8e-07 W=4.4e-07 $X=-7990 $Y=-6960 $D=4
M491 VDD 197 204 VDD PM L=1.8e-07 W=8.8e-07 $X=-7800 $Y=-30500 $D=4
M492 VDD 57 207 VDD PM L=1.8e-07 W=8.8e-07 $X=-7650 $Y=-56400 $D=4
M493 VDD 58 210 VDD PM L=1.8e-07 W=8.8e-07 $X=-7650 $Y=5550 $D=4
M494 VDD 33 462 VDD PM L=1.8e-07 W=8.8e-07 $X=-7530 $Y=-46250 $D=4
M495 VDD 34 463 VDD PM L=1.8e-07 W=8.8e-07 $X=-7530 $Y=-4600 $D=4
M496 198 35 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-7080 $Y=-19910 $D=4
M497 464 57 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6930 $Y=-56400 $D=4
M498 465 58 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-6930 $Y=5550 $D=4
M499 466 59 464 VDD PM L=1.8e-07 W=8.8e-07 $X=-6500 $Y=-56400 $D=4
M500 467 60 465 VDD PM L=1.8e-07 W=8.8e-07 $X=-6500 $Y=5550 $D=4
M501 240 46 466 VDD PM L=1.8e-07 W=8.8e-07 $X=-6070 $Y=-56400 $D=4
M502 241 47 467 VDD PM L=1.8e-07 W=8.8e-07 $X=-6070 $Y=5550 $D=4
M503 227 75 36 VDD PM L=1.8e-07 W=4.4e-07 $X=-5940 $Y=-43450 $D=4
M504 228 76 37 VDD PM L=1.8e-07 W=4.4e-07 $X=-5940 $Y=-6960 $D=4
M505 225 71 36 VDD PM L=1.8e-07 W=4.4e-07 $X=-5890 $Y=-32860 $D=4
M506 226 72 37 VDD PM L=1.8e-07 W=4.4e-07 $X=-5890 $Y=-17550 $D=4
M507 233 215 240 VDD PM L=1.8e-07 W=8.8e-07 $X=-5350 $Y=-56400 $D=4
M508 236 216 241 VDD PM L=1.8e-07 W=8.8e-07 $X=-5350 $Y=5550 $D=4
M509 VDD 46 233 VDD PM L=1.8e-07 W=8.8e-07 $X=-4630 $Y=-56400 $D=4
M510 VDD 47 236 VDD PM L=1.8e-07 W=8.8e-07 $X=-4630 $Y=5550 $D=4
M511 229 198 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-4420 $Y=-19910 $D=4
M512 230 75 48 VDD PM L=1.8e-07 W=4.4e-07 $X=-3990 $Y=-43450 $D=4
M513 231 35 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-3990 $Y=-30500 $D=4
M514 232 76 49 VDD PM L=1.8e-07 W=4.4e-07 $X=-3990 $Y=-6960 $D=4
M515 237 71 48 VDD PM L=1.8e-07 W=4.4e-07 $X=-3950 $Y=-32860 $D=4
M516 233 59 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-3910 $Y=-56400 $D=4
M517 236 60 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-3910 $Y=5550 $D=4
M518 468 35 229 VDD PM L=1.8e-07 W=8.8e-07 $X=-3660 $Y=-20350 $D=4
M519 VDD 261 63 VDD PM L=1.8e-07 W=8.8e-07 $X=-3610 $Y=-46250 $D=4
M520 VDD 262 64 VDD PM L=1.8e-07 W=8.8e-07 $X=-3610 $Y=-4600 $D=4
M521 GND B0 50 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-69640 $D=4
M522 GND B0 101 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-65160 $D=4
M523 GND B0 115 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-63020 $D=4
M524 GND B0 129 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=-58540 $D=4
M525 GND X0 130 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=8350 $D=4
M526 GND X0 116 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=12830 $D=4
M527 GND X0 102 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=14970 $D=4
M528 GND X0 51 VDD PM L=1.8e-07 W=2.2e-07 $X=-3300 $Y=19450 $D=4
M529 VDD 52 468 VDD PM L=1.8e-07 W=8.8e-07 $X=-3230 $Y=-20350 $D=4
M530 VDD 57 233 VDD PM L=1.8e-07 W=8.8e-07 $X=-3190 $Y=-56400 $D=4
M531 VDD 225 237 VDD PM L=1.8e-07 W=8.8e-07 $X=-3190 $Y=-33300 $D=4
M532 VDD 226 238 VDD PM L=1.8e-07 W=8.8e-07 $X=-3190 $Y=-17550 $D=4
M533 VDD 58 236 VDD PM L=1.8e-07 W=8.8e-07 $X=-3190 $Y=5550 $D=4
M534 66 240 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-2470 $Y=-56400 $D=4
M535 227 55 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=-43450 $D=4
M536 469 63 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-2470 $Y=-33300 $D=4
M537 228 56 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-2470 $Y=-6960 $D=4
M538 67 241 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-2470 $Y=5550 $D=4
M539 226 56 470 VDD PM L=1.8e-07 W=8.8e-07 $X=-2040 $Y=-17550 $D=4
M540 VDD 69 246 VDD PM L=1.8e-07 W=8.8e-07 $X=-1670 $Y=-46250 $D=4
M541 VDD 70 247 VDD PM L=1.8e-07 W=8.8e-07 $X=-1670 $Y=-4600 $D=4
M542 243 242 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-1330 $Y=-30500 $D=4
M543 471 69 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-950 $Y=-46250 $D=4
M544 472 70 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-950 $Y=-4600 $D=4
M545 O6 62 243 VDD PM L=1.8e-07 W=4.4e-07 $X=-570 $Y=-30500 $D=4
M546 O6 65 244 VDD PM L=1.8e-07 W=4.4e-07 $X=-530 $Y=-19910 $D=4
M547 261 73 471 VDD PM L=1.8e-07 W=8.8e-07 $X=-520 $Y=-46250 $D=4
M548 262 74 472 VDD PM L=1.8e-07 W=8.8e-07 $X=-520 $Y=-4600 $D=4
M549 VDD 64 252 VDD PM L=1.8e-07 W=8.8e-07 $X=-100 $Y=-17550 $D=4
M550 249 227 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=190 $Y=-43450 $D=4
M551 250 228 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=190 $Y=-6960 $D=4
M552 246 66 261 VDD PM L=1.8e-07 W=8.8e-07 $X=200 $Y=-46250 $D=4
M553 247 67 262 VDD PM L=1.8e-07 W=8.8e-07 $X=200 $Y=-4600 $D=4
M554 253 53 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=270 $Y=-56400 $D=4
M555 254 54 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=270 $Y=5990 $D=4
M556 251 55 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=620 $Y=-33300 $D=4
M557 252 56 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=620 $Y=-17550 $D=4
M558 VDD 73 246 VDD PM L=1.8e-07 W=8.8e-07 $X=920 $Y=-46250 $D=4
M559 VDD 74 247 VDD PM L=1.8e-07 W=8.8e-07 $X=920 $Y=-4600 $D=4
M560 260 88 62 VDD PM L=1.8e-07 W=4.4e-07 $X=1520 $Y=-19910 $D=4
M561 259 85 62 VDD PM L=1.8e-07 W=4.4e-07 $X=1570 $Y=-30500 $D=4
M562 473 73 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=1640 $Y=-46250 $D=4
M563 474 74 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=1640 $Y=-4600 $D=4
M564 475 69 473 VDD PM L=1.8e-07 W=8.8e-07 $X=2070 $Y=-46250 $D=4
M565 476 70 474 VDD PM L=1.8e-07 W=8.8e-07 $X=2070 $Y=-4600 $D=4
M566 277 66 475 VDD PM L=1.8e-07 W=8.8e-07 $X=2500 $Y=-46250 $D=4
M567 278 67 476 VDD PM L=1.8e-07 W=8.8e-07 $X=2500 $Y=-4600 $D=4
M568 263 253 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=2930 $Y=-56400 $D=4
M569 264 254 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=2930 $Y=5990 $D=4
M570 274 261 277 VDD PM L=1.8e-07 W=8.8e-07 $X=3220 $Y=-46250 $D=4
M571 275 262 278 VDD PM L=1.8e-07 W=8.8e-07 $X=3220 $Y=-4600 $D=4
M572 265 257 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=3280 $Y=-33300 $D=4
M573 266 258 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=3280 $Y=-17550 $D=4
M574 267 249 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=3320 $Y=-43450 $D=4
M575 268 250 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=3320 $Y=-7400 $D=4
M576 269 88 65 VDD PM L=1.8e-07 W=4.4e-07 $X=3470 $Y=-19910 $D=4
M577 VDD 66 274 VDD PM L=1.8e-07 W=8.8e-07 $X=3940 $Y=-46250 $D=4
M578 VDD 67 275 VDD PM L=1.8e-07 W=8.8e-07 $X=3940 $Y=-4600 $D=4
M579 78 71 265 VDD PM L=1.8e-07 W=4.4e-07 $X=4040 $Y=-32860 $D=4
M580 68 72 266 VDD PM L=1.8e-07 W=4.4e-07 $X=4040 $Y=-17550 $D=4
M581 78 75 267 VDD PM L=1.8e-07 W=4.4e-07 $X=4080 $Y=-43450 $D=4
M582 68 76 268 VDD PM L=1.8e-07 W=4.4e-07 $X=4080 $Y=-6960 $D=4
M583 VDD 259 270 VDD PM L=1.8e-07 W=8.8e-07 $X=4270 $Y=-30500 $D=4
M584 274 69 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=4660 $Y=-46250 $D=4
M585 275 70 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=4660 $Y=-4600 $D=4
M586 260 68 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=4990 $Y=-19910 $D=4
M587 VDD 73 274 VDD PM L=1.8e-07 W=8.8e-07 $X=5380 $Y=-46250 $D=4
M588 VDD 74 275 VDD PM L=1.8e-07 W=8.8e-07 $X=5380 $Y=-4600 $D=4
M589 VDD 78 260 VDD PM L=1.8e-07 W=4.4e-07 $X=5710 $Y=-19910 $D=4
M590 80 277 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=6100 $Y=-46250 $D=4
M591 81 278 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=6100 $Y=-4600 $D=4
M592 279 283 71 VDD PM L=1.8e-07 W=4.4e-07 $X=6180 $Y=-32860 $D=4
M593 VDD 78 289 VDD PM L=1.8e-07 W=8.8e-07 $X=7360 $Y=-30500 $D=4
M594 287 260 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=7650 $Y=-19910 $D=4
M595 VDD 317 82 VDD PM L=1.8e-07 W=8.8e-07 $X=8040 $Y=-46250 $D=4
M596 VDD 318 83 VDD PM L=1.8e-07 W=8.8e-07 $X=8040 $Y=-4600 $D=4
M597 288 285 75 VDD PM L=1.8e-07 W=4.4e-07 $X=8080 $Y=-43450 $D=4
M598 289 68 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=8080 $Y=-30500 $D=4
M599 290 286 76 VDD PM L=1.8e-07 W=4.4e-07 $X=8080 $Y=-6960 $D=4
M600 291 283 75 VDD PM L=1.8e-07 W=4.4e-07 $X=8120 $Y=-32860 $D=4
M601 292 284 76 VDD PM L=1.8e-07 W=4.4e-07 $X=8120 $Y=-17550 $D=4
M602 294 259 289 VDD PM L=1.8e-07 W=8.8e-07 $X=8800 $Y=-30500 $D=4
M603 295 77 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=8840 $Y=-56400 $D=4
M604 296 79 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=8840 $Y=5990 $D=4
M605 VDD 279 291 VDD PM L=1.8e-07 W=8.8e-07 $X=8880 $Y=-33300 $D=4
M606 VDD 280 292 VDD PM L=1.8e-07 W=8.8e-07 $X=8880 $Y=-17550 $D=4
M607 281 80 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=9600 $Y=-43450 $D=4
M608 477 83 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=9600 $Y=-17550 $D=4
M609 282 81 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=9600 $Y=-6960 $D=4
M610 VDD 91 302 VDD PM L=1.8e-07 W=8.8e-07 $X=9980 $Y=-46250 $D=4
M611 VDD 92 303 VDD PM L=1.8e-07 W=8.8e-07 $X=9980 $Y=-4600 $D=4
M612 478 91 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10700 $Y=-46250 $D=4
M613 479 92 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10700 $Y=-4600 $D=4
M614 297 294 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10740 $Y=-30500 $D=4
M615 298 287 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10780 $Y=-20350 $D=4
M616 317 93 478 VDD PM L=1.8e-07 W=8.8e-07 $X=11130 $Y=-46250 $D=4
M617 318 94 479 VDD PM L=1.8e-07 W=8.8e-07 $X=11130 $Y=-4600 $D=4
M618 299 295 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=11500 $Y=-56400 $D=4
M619 O5 85 297 VDD PM L=1.8e-07 W=4.4e-07 $X=11500 $Y=-30500 $D=4
M620 300 296 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=11500 $Y=5990 $D=4
M621 O5 88 298 VDD PM L=1.8e-07 W=4.4e-07 $X=11540 $Y=-19910 $D=4
M622 302 89 317 VDD PM L=1.8e-07 W=8.8e-07 $X=11850 $Y=-46250 $D=4
M623 303 90 318 VDD PM L=1.8e-07 W=8.8e-07 $X=11850 $Y=-4600 $D=4
M624 305 281 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=12260 $Y=-43450 $D=4
M625 306 282 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=12260 $Y=-6960 $D=4
M626 VDD 93 302 VDD PM L=1.8e-07 W=8.8e-07 $X=12570 $Y=-46250 $D=4
M627 VDD 94 303 VDD PM L=1.8e-07 W=8.8e-07 $X=12570 $Y=-4600 $D=4
M628 309 80 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=12690 $Y=-33300 $D=4
M629 310 81 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=12690 $Y=-17550 $D=4
M630 480 93 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=13290 $Y=-46250 $D=4
M631 481 94 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=13290 $Y=-4600 $D=4
M632 313 279 309 VDD PM L=1.8e-07 W=8.8e-07 $X=13410 $Y=-33300 $D=4
M633 316 109 85 VDD PM L=1.8e-07 W=4.4e-07 $X=13590 $Y=-19910 $D=4
M634 482 91 480 VDD PM L=1.8e-07 W=8.8e-07 $X=13720 $Y=-46250 $D=4
M635 483 92 481 VDD PM L=1.8e-07 W=8.8e-07 $X=13720 $Y=-4600 $D=4
M636 329 89 482 VDD PM L=1.8e-07 W=8.8e-07 $X=14150 $Y=-46250 $D=4
M637 330 90 483 VDD PM L=1.8e-07 W=8.8e-07 $X=14150 $Y=-4600 $D=4
M638 326 317 329 VDD PM L=1.8e-07 W=8.8e-07 $X=14870 $Y=-46250 $D=4
M639 327 318 330 VDD PM L=1.8e-07 W=8.8e-07 $X=14870 $Y=-4600 $D=4
M640 320 314 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=15350 $Y=-17550 $D=4
M641 323 109 88 VDD PM L=1.8e-07 W=4.4e-07 $X=15540 $Y=-19910 $D=4
M642 324 106 88 VDD PM L=1.8e-07 W=4.4e-07 $X=15580 $Y=-30500 $D=4
M643 VDD 89 326 VDD PM L=1.8e-07 W=8.8e-07 $X=15590 $Y=-46250 $D=4
M644 VDD 90 327 VDD PM L=1.8e-07 W=8.8e-07 $X=15590 $Y=-4600 $D=4
M645 98 283 319 VDD PM L=1.8e-07 W=4.4e-07 $X=16110 $Y=-32860 $D=4
M646 95 284 320 VDD PM L=1.8e-07 W=4.4e-07 $X=16110 $Y=-17550 $D=4
M647 98 285 321 VDD PM L=1.8e-07 W=4.4e-07 $X=16150 $Y=-43450 $D=4
M648 95 286 322 VDD PM L=1.8e-07 W=4.4e-07 $X=16150 $Y=-6960 $D=4
M649 326 91 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=16310 $Y=-46250 $D=4
M650 327 92 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=16310 $Y=-4600 $D=4
M651 VDD 315 324 VDD PM L=1.8e-07 W=8.8e-07 $X=16340 $Y=-30500 $D=4
M652 VDD 347 89 VDD PM L=1.8e-07 W=8.8e-07 $X=16610 $Y=-56400 $D=4
M653 VDD 348 90 VDD PM L=1.8e-07 W=8.8e-07 $X=16610 $Y=5550 $D=4
M654 VDD 93 326 VDD PM L=1.8e-07 W=8.8e-07 $X=17030 $Y=-46250 $D=4
M655 VDD 94 327 VDD PM L=1.8e-07 W=8.8e-07 $X=17030 $Y=-4600 $D=4
M656 316 95 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17060 $Y=-19910 $D=4
M657 99 329 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=17750 $Y=-46250 $D=4
M658 100 330 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=17750 $Y=-4600 $D=4
M659 VDD 104 333 VDD PM L=1.8e-07 W=8.8e-07 $X=18550 $Y=-56400 $D=4
M660 VDD 105 336 VDD PM L=1.8e-07 W=8.8e-07 $X=18550 $Y=5550 $D=4
M661 283 96 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18890 $Y=-43450 $D=4
M662 284 97 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18890 $Y=-6960 $D=4
M663 484 104 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=19270 $Y=-56400 $D=4
M664 485 105 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=19270 $Y=5550 $D=4
M665 VDD 99 283 VDD PM L=1.8e-07 W=4.4e-07 $X=19610 $Y=-43450 $D=4
M666 VDD 100 284 VDD PM L=1.8e-07 W=4.4e-07 $X=19610 $Y=-6960 $D=4
M667 347 31 484 VDD PM L=1.8e-07 W=8.8e-07 $X=19700 $Y=-56400 $D=4
M668 348 32 485 VDD PM L=1.8e-07 W=8.8e-07 $X=19700 $Y=5550 $D=4
M669 331 316 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=19720 $Y=-19910 $D=4
M670 332 95 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=20150 $Y=-30500 $D=4
M671 333 101 347 VDD PM L=1.8e-07 W=8.8e-07 $X=20420 $Y=-56400 $D=4
M672 336 102 348 VDD PM L=1.8e-07 W=8.8e-07 $X=20420 $Y=5550 $D=4
M673 339 110 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20490 $Y=-45810 $D=4
M674 340 111 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20490 $Y=-4600 $D=4
M675 VDD 31 333 VDD PM L=1.8e-07 W=8.8e-07 $X=21140 $Y=-56400 $D=4
M676 VDD 32 336 VDD PM L=1.8e-07 W=8.8e-07 $X=21140 $Y=5550 $D=4
M677 341 283 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=21550 $Y=-43450 $D=4
M678 342 284 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=21550 $Y=-6960 $D=4
M679 486 31 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=21860 $Y=-56400 $D=4
M680 487 32 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=21860 $Y=5550 $D=4
M681 488 104 486 VDD PM L=1.8e-07 W=8.8e-07 $X=22290 $Y=-56400 $D=4
M682 489 105 487 VDD PM L=1.8e-07 W=8.8e-07 $X=22290 $Y=5550 $D=4
M683 357 101 488 VDD PM L=1.8e-07 W=8.8e-07 $X=22720 $Y=-56400 $D=4
M684 358 102 489 VDD PM L=1.8e-07 W=8.8e-07 $X=22720 $Y=5550 $D=4
M685 349 339 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23150 $Y=-45810 $D=4
M686 350 340 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23150 $Y=-4600 $D=4
M687 353 347 357 VDD PM L=1.8e-07 W=8.8e-07 $X=23440 $Y=-56400 $D=4
M688 356 348 358 VDD PM L=1.8e-07 W=8.8e-07 $X=23440 $Y=5550 $D=4
M689 O4 106 345 VDD PM L=1.8e-07 W=4.4e-07 $X=23570 $Y=-30500 $D=4
M690 O4 109 346 VDD PM L=1.8e-07 W=4.4e-07 $X=23610 $Y=-19910 $D=4
M691 VDD 101 353 VDD PM L=1.8e-07 W=8.8e-07 $X=24160 $Y=-56400 $D=4
M692 VDD 102 356 VDD PM L=1.8e-07 W=8.8e-07 $X=24160 $Y=5550 $D=4
M693 117 341 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=24680 $Y=-43450 $D=4
M694 114 342 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=24680 $Y=-6960 $D=4
M695 353 104 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=24880 $Y=-56400 $D=4
M696 356 105 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=24880 $Y=5550 $D=4
M697 VDD 31 353 VDD PM L=1.8e-07 W=8.8e-07 $X=25600 $Y=-56400 $D=4
M698 VDD 32 356 VDD PM L=1.8e-07 W=8.8e-07 $X=25600 $Y=5550 $D=4
M699 107 357 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=26320 $Y=-56400 $D=4
M700 108 358 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=26320 $Y=5550 $D=4
M701 361 120 109 VDD PM L=1.8e-07 W=4.4e-07 $X=27610 $Y=-19910 $D=4
M702 VDD 359 362 VDD PM L=1.8e-07 W=8.8e-07 $X=28410 $Y=-30500 $D=4
M703 363 112 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29060 $Y=-56400 $D=4
M704 364 113 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29060 $Y=5990 $D=4
M705 360 114 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29130 $Y=-19910 $D=4
M706 365 363 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31720 $Y=-56400 $D=4
M707 366 364 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31720 $Y=5990 $D=4
M708 367 360 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31790 $Y=-19910 $D=4
M709 368 114 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=32220 $Y=-30500 $D=4
M710 O3 119 373 VDD PM L=1.8e-07 W=4.4e-07 $X=35640 $Y=-30500 $D=4
M711 O3 120 374 VDD PM L=1.8e-07 W=4.4e-07 $X=35680 $Y=-19910 $D=4
M712 377 125 120 VDD PM L=1.8e-07 W=4.4e-07 $X=39680 $Y=-19910 $D=4
M713 VDD 375 378 VDD PM L=1.8e-07 W=8.8e-07 $X=40480 $Y=-30500 $D=4
M714 376 121 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=41200 $Y=-19910 $D=4
M715 379 376 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=43860 $Y=-19910 $D=4
M716 380 121 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44290 $Y=-30500 $D=4
M717 O2 124 383 VDD PM L=1.8e-07 W=4.4e-07 $X=47710 $Y=-30500 $D=4
M718 O2 125 384 VDD PM L=1.8e-07 W=4.4e-07 $X=47750 $Y=-19910 $D=4
M719 389 388 125 VDD PM L=1.8e-07 W=4.4e-07 $X=51750 $Y=-19910 $D=4
M720 VDD 385 390 VDD PM L=1.8e-07 W=8.8e-07 $X=52550 $Y=-30500 $D=4
M721 386 126 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=53270 $Y=-19910 $D=4
M722 391 386 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=55930 $Y=-19910 $D=4
M723 392 126 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=56360 $Y=-30500 $D=4
M724 O1 387 395 VDD PM L=1.8e-07 W=4.4e-07 $X=59780 $Y=-30500 $D=4
M725 O1 388 396 VDD PM L=1.8e-07 W=4.4e-07 $X=59820 $Y=-19910 $D=4
M726 387 129 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=62560 $Y=-19910 $D=4
M727 397 387 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=65220 $Y=-19910 $D=4
X728 VDD 3 19 15 p18_CDNS_672684331922 $T=-20670 -43010 1 0 $X=-21580 $Y=-44800
X729 VDD 4 12 16 p18_CDNS_672684331922 $T=-20670 -6960 0 0 $X=-21580 $Y=-7390
X730 VDD 132 O8 29 p18_CDNS_672684331922 $T=-20450 -30060 0 180 $X=-21540 $Y=-31850
X731 VDD 13 147 48 p18_CDNS_672684331922 $T=-18010 -43010 1 0 $X=-18920 $Y=-44800
X732 VDD 14 148 49 p18_CDNS_672684331922 $T=-18010 -6960 0 0 $X=-18920 $Y=-7390
X733 VDD 145 13 36 p18_CDNS_672684331922 $T=-17780 -32860 1 180 $X=-18870 $Y=-33290
X734 VDD 146 14 37 p18_CDNS_672684331922 $T=-17780 -17110 0 180 $X=-18870 $Y=-18900
X735 VDD 164 16 37 p18_CDNS_672684331922 $T=-15840 -17110 0 180 $X=-16930 $Y=-18900
X736 VDD VDD 33 149 p18_CDNS_672684331922 $T=-14160 -55960 1 0 $X=-15070 $Y=-57750
X737 VDD VDD 20 150 p18_CDNS_672684331922 $T=-14160 -45810 0 0 $X=-15070 $Y=-46240
X738 VDD VDD 21 151 p18_CDNS_672684331922 $T=-14160 -4160 1 0 $X=-15070 $Y=-5950
X739 VDD VDD 34 152 p18_CDNS_672684331922 $T=-14160 5990 0 0 $X=-15070 $Y=5560
X740 VDD 24 VDD 185 p18_CDNS_672684331922 $T=-12100 -45810 0 0 $X=-13010 $Y=-46240
X741 VDD 25 VDD 186 p18_CDNS_672684331922 $T=-12100 -4160 1 0 $X=-13010 $Y=-5950
X742 VDD 204 30 62 p18_CDNS_672684331922 $T=-8380 -30060 0 180 $X=-9470 $Y=-31850
X743 VDD 198 VDD 52 p18_CDNS_672684331922 $T=-6360 -19910 0 0 $X=-7270 $Y=-20340
X744 VDD VDD 55 205 p18_CDNS_672684331922 $T=-5590 -45810 0 0 $X=-6500 $Y=-46240
X745 VDD VDD 56 206 p18_CDNS_672684331922 $T=-5590 -4160 1 0 $X=-6500 $Y=-5950
X746 VDD 238 49 72 p18_CDNS_672684331922 $T=-3770 -17110 0 180 $X=-4860 $Y=-18900
X747 VDD 227 VDD 63 p18_CDNS_672684331922 $T=-1750 -43010 1 0 $X=-2660 $Y=-44800
X748 VDD 228 VDD 64 p18_CDNS_672684331922 $T=-1750 -6960 0 0 $X=-2660 $Y=-7390
X749 VDD 270 65 85 p18_CDNS_672684331922 $T=3690 -30060 0 180 $X=2600 $Y=-31850
X750 VDD VDD 93 263 p18_CDNS_672684331922 $T=6060 -55960 1 0 $X=5150 $Y=-57750
X751 VDD VDD 94 264 p18_CDNS_672684331922 $T=6060 5990 0 0 $X=5150 $Y=5560
X752 VDD 71 281 285 p18_CDNS_672684331922 $T=6130 -43010 1 0 $X=5220 $Y=-44800
X753 VDD 72 282 286 p18_CDNS_672684331922 $T=6130 -6960 0 0 $X=5220 $Y=-7390
X754 VDD 280 72 284 p18_CDNS_672684331922 $T=6360 -17110 0 180 $X=5270 $Y=-18900
X755 VDD 281 VDD 82 p18_CDNS_672684331922 $T=10320 -43010 1 0 $X=9410 $Y=-44800
X756 VDD 282 VDD 83 p18_CDNS_672684331922 $T=10320 -6960 0 0 $X=9410 $Y=-7390
X757 VDD 315 85 106 p18_CDNS_672684331922 $T=13820 -30060 0 180 $X=12730 $Y=-31850
X758 VDD VDD 91 299 p18_CDNS_672684331922 $T=14630 -55960 1 0 $X=13720 $Y=-57750
X759 VDD VDD 92 300 p18_CDNS_672684331922 $T=14630 5990 0 0 $X=13720 $Y=5560
X760 VDD 316 VDD 98 p18_CDNS_672684331922 $T=17780 -19910 0 0 $X=16870 $Y=-20340
X761 VDD 285 VDD 283 p18_CDNS_672684331922 $T=18170 -43010 1 0 $X=17260 $Y=-44800
X762 VDD 286 VDD 284 p18_CDNS_672684331922 $T=18170 -6960 0 0 $X=17260 $Y=-7390
X763 VDD 106 360 120 p18_CDNS_672684331922 $T=25660 -19910 0 0 $X=24750 $Y=-20340
X764 VDD 359 106 119 p18_CDNS_672684331922 $T=25890 -30060 0 180 $X=24800 $Y=-31850
X765 VDD VDD 122 349 p18_CDNS_672684331922 $T=26280 -45810 0 0 $X=25370 $Y=-46240
X766 VDD VDD 121 350 p18_CDNS_672684331922 $T=26280 -4160 1 0 $X=25370 $Y=-5950
X767 VDD 362 109 119 p18_CDNS_672684331922 $T=27830 -30060 0 180 $X=26740 $Y=-31850
X768 VDD 360 VDD 117 p18_CDNS_672684331922 $T=29850 -19910 0 0 $X=28940 $Y=-20340
X769 VDD VDD 127 365 p18_CDNS_672684331922 $T=34850 -55960 1 0 $X=33940 $Y=-57750
X770 VDD VDD 126 366 p18_CDNS_672684331922 $T=34850 5990 0 0 $X=33940 $Y=5560
X771 VDD 119 376 125 p18_CDNS_672684331922 $T=37730 -19910 0 0 $X=36820 $Y=-20340
X772 VDD 375 119 124 p18_CDNS_672684331922 $T=37960 -30060 0 180 $X=36870 $Y=-31850
X773 VDD 378 120 124 p18_CDNS_672684331922 $T=39900 -30060 0 180 $X=38810 $Y=-31850
X774 VDD 376 VDD 122 p18_CDNS_672684331922 $T=41920 -19910 0 0 $X=41010 $Y=-20340
X775 VDD 124 386 388 p18_CDNS_672684331922 $T=49800 -19910 0 0 $X=48890 $Y=-20340
X776 VDD 385 124 387 p18_CDNS_672684331922 $T=50030 -30060 0 180 $X=48940 $Y=-31850
X777 VDD 390 125 387 p18_CDNS_672684331922 $T=51970 -30060 0 180 $X=50880 $Y=-31850
X778 VDD 386 VDD 127 p18_CDNS_672684331922 $T=53990 -19910 0 0 $X=53080 $Y=-20340
X779 VDD VDD O0 397 p18_CDNS_672684331922 $T=68350 -19910 0 0 $X=67440 $Y=-20340
X780 VDD VDD 19 452 p18_CDNS_672684331923 $T=-19150 -29620 1 0 $X=-20060 $Y=-31850
X781 VDD 150 6 453 p18_CDNS_672684331923 $T=-16530 -46250 0 0 $X=-17440 $Y=-46680
X782 VDD 151 7 454 p18_CDNS_672684331923 $T=-16530 -3720 1 0 $X=-17440 $Y=-5950
X783 VDD VDD 24 457 p18_CDNS_672684331923 $T=-14540 -33300 0 0 $X=-15450 $Y=-33730
X784 VDD 179 20 458 p18_CDNS_672684331923 $T=-11120 -42570 1 0 $X=-12030 $Y=-44800
X785 VDD 180 21 459 p18_CDNS_672684331923 $T=-11120 -7400 0 0 $X=-12030 $Y=-7830
X786 VDD 205 27 462 p18_CDNS_672684331923 $T=-7960 -46250 0 0 $X=-8870 $Y=-46680
X787 VDD 206 28 463 p18_CDNS_672684331923 $T=-7960 -3720 1 0 $X=-8870 $Y=-5950
X788 VDD VDD 64 470 p18_CDNS_672684331923 $T=-2470 -16670 1 0 $X=-3380 $Y=-18900
X789 VDD VDD 19 455 p18_CDNS_672684331928 $T=-15300 -20350 0 0 $X=-15855 $Y=-20780
X790 VDD 146 21 456 p18_CDNS_672684331928 $T=-14110 -16670 1 0 $X=-14665 $Y=-18900
X791 VDD 225 55 469 p18_CDNS_672684331928 $T=-2040 -33300 0 0 $X=-2595 $Y=-33730
X792 VDD 280 81 477 p18_CDNS_672684331928 $T=10030 -16670 1 0 $X=9475 $Y=-18900
X793 VDD 149 VDD 8 22 ICV_1 $T=-16530 -55520 1 0 $X=-17440 $Y=-57750
X794 VDD 152 VDD 9 23 ICV_1 $T=-16530 5550 0 0 $X=-17440 $Y=5120
X795 VDD VDD 197 52 35 ICV_1 $T=-7080 -29620 1 0 $X=-7990 $Y=-31850
X796 VDD 249 VDD 55 63 ICV_1 $T=950 -42570 1 0 $X=40 $Y=-44800
X797 VDD 250 VDD 56 64 ICV_1 $T=950 -7400 0 0 $X=40 $Y=-7830
X798 VDD 263 VDD 53 50 ICV_1 $T=3690 -55520 1 0 $X=2780 $Y=-57750
X799 VDD 264 VDD 54 51 ICV_1 $T=3690 5550 0 0 $X=2780 $Y=5120
X800 VDD VDD 259 78 68 ICV_1 $T=4990 -29620 1 0 $X=4080 $Y=-31850
X801 VDD 287 VDD 68 78 ICV_1 $T=8410 -20350 0 0 $X=7500 $Y=-20780
X802 VDD VDD 279 82 80 ICV_1 $T=9600 -33300 0 0 $X=8690 $Y=-33730
X803 VDD 299 VDD 77 86 ICV_1 $T=12260 -55520 1 0 $X=11350 $Y=-57750
X804 VDD 300 VDD 79 87 ICV_1 $T=12260 5550 0 0 $X=11350 $Y=5120
X805 VDD 305 VDD 80 82 ICV_1 $T=13020 -42570 1 0 $X=12110 $Y=-44800
X806 VDD 306 VDD 81 83 ICV_1 $T=13020 -7400 0 0 $X=12110 $Y=-7830
X807 VDD VDD 315 98 95 ICV_1 $T=17060 -29620 1 0 $X=16150 $Y=-31850
X808 VDD 331 VDD 95 98 ICV_1 $T=20480 -20350 0 0 $X=19570 $Y=-20780
X809 VDD 341 VDD 96 99 ICV_1 $T=22310 -42570 1 0 $X=21400 $Y=-44800
X810 VDD 342 VDD 97 100 ICV_1 $T=22310 -7400 0 0 $X=21400 $Y=-7830
X811 VDD 349 VDD 110 107 ICV_1 $T=23910 -46250 0 0 $X=23000 $Y=-46680
X812 VDD 350 VDD 111 108 ICV_1 $T=23910 -3720 1 0 $X=23000 $Y=-5950
X813 VDD VDD 359 117 114 ICV_1 $T=29130 -29620 1 0 $X=28220 $Y=-31850
X814 VDD 365 VDD 112 115 ICV_1 $T=32480 -55520 1 0 $X=31570 $Y=-57750
X815 VDD 366 VDD 113 116 ICV_1 $T=32480 5550 0 0 $X=31570 $Y=5120
X816 VDD 367 VDD 114 117 ICV_1 $T=32550 -20350 0 0 $X=31640 $Y=-20780
X817 VDD VDD 375 122 121 ICV_1 $T=41200 -29620 1 0 $X=40290 $Y=-31850
X818 VDD 379 VDD 121 122 ICV_1 $T=44620 -20350 0 0 $X=43710 $Y=-20780
X819 VDD VDD 385 127 126 ICV_1 $T=53270 -29620 1 0 $X=52360 $Y=-31850
X820 VDD 391 VDD 126 127 ICV_1 $T=56690 -20350 0 0 $X=55780 $Y=-20780
X821 VDD 397 VDD 129 130 ICV_1 $T=65980 -20350 0 0 $X=65070 $Y=-20780
X822 GND 3 19 13 n18_CDNS_672684331926 $T=-20670 -39565 1 0 $X=-21330 $Y=-40355
X823 GND 131 O8 29 n18_CDNS_672684331926 $T=-20490 -23355 1 180 $X=-21330 $Y=-25375
X824 GND 4 12 14 n18_CDNS_672684331926 $T=-20670 -10405 0 0 $X=-21330 $Y=-12425
X825 GND 98 321 283 n18_CDNS_672684331926 $T=16330 -39565 0 180 $X=15490 $Y=-40355
X826 GND 95 322 284 n18_CDNS_672684331926 $T=16330 -10405 1 180 $X=15490 $Y=-12425
X827 GND O1 396 387 n18_CDNS_672684331926 $T=60000 -23355 1 180 $X=59160 $Y=-25375
X828 GND 141 149 156 8 22 ICV_2 $T=-19950 -52515 1 0 $X=-20610 $Y=-53305
X829 GND 10 150 157 6 17 ICV_2 $T=-19950 -49255 0 0 $X=-20610 $Y=-51275
X830 GND 11 151 158 7 18 ICV_2 $T=-19950 -715 1 0 $X=-20610 $Y=-1505
X831 GND 142 152 159 9 23 ICV_2 $T=-19950 2545 0 0 $X=-20610 $Y=525
X832 GND 185 205 211 27 33 ICV_2 $T=-11380 -49255 0 0 $X=-12040 $Y=-51275
X833 GND 186 206 212 28 34 ICV_2 $T=-11380 -715 1 0 $X=-12040 $Y=-1505
X834 GND 253 263 271 53 50 ICV_2 $T=270 -52515 1 0 $X=-390 $Y=-53305
X835 GND 254 264 272 54 51 ICV_2 $T=270 2545 0 0 $X=-390 $Y=525
X836 GND 295 299 307 77 86 ICV_2 $T=8840 -52515 1 0 $X=8180 $Y=-53305
X837 GND 296 300 308 79 87 ICV_2 $T=8840 2545 0 0 $X=8180 $Y=525
X838 GND 283 341 343 96 99 ICV_2 $T=18890 -39565 1 0 $X=18230 $Y=-40355
X839 GND 284 342 344 97 100 ICV_2 $T=18890 -10405 0 0 $X=18230 $Y=-12425
X840 GND 339 349 351 110 107 ICV_2 $T=20490 -49255 0 0 $X=19830 $Y=-51275
X841 GND 340 350 352 111 108 ICV_2 $T=20490 -715 1 0 $X=19830 $Y=-1505
X842 GND 363 365 369 112 115 ICV_2 $T=29060 -52515 1 0 $X=28400 $Y=-53305
X843 GND 364 366 370 113 116 ICV_2 $T=29060 2545 0 0 $X=28400 $Y=525
X844 GND 387 397 398 129 130 ICV_2 $T=62560 -23355 0 0 $X=61900 $Y=-25375
X845 VDD 6 141 22 ICV_3 $T=-20670 -55960 1 0 $X=-21580 $Y=-57750
X846 VDD 3 10 17 ICV_3 $T=-20670 -45810 0 0 $X=-21580 $Y=-46240
X847 VDD 4 11 18 ICV_3 $T=-20670 -4160 1 0 $X=-21580 $Y=-5950
X848 VDD 7 142 23 ICV_3 $T=-20670 5990 0 0 $X=-21580 $Y=5560
X849 VDD 73 253 50 ICV_3 $T=-450 -55960 1 0 $X=-1360 $Y=-57750
X850 VDD 74 254 51 ICV_3 $T=-450 5990 0 0 $X=-1360 $Y=5560
X851 VDD 69 295 86 ICV_3 $T=8120 -55960 1 0 $X=7210 $Y=-57750
X852 VDD 70 296 87 ICV_3 $T=8120 5990 0 0 $X=7210 $Y=5560
X853 VDD 96 339 107 ICV_3 $T=19770 -45810 0 0 $X=18860 $Y=-46240
X854 VDD 97 340 108 ICV_3 $T=19770 -4160 1 0 $X=18860 $Y=-5950
X855 VDD 110 363 115 ICV_3 $T=28340 -55960 1 0 $X=27430 $Y=-57750
X856 VDD 111 364 116 ICV_3 $T=28340 5990 0 0 $X=27430 $Y=5560
X857 VDD 388 387 130 ICV_3 $T=61840 -19910 0 0 $X=60930 $Y=-20340
X858 VDD 131 VDD 144 p18_CDNS_6726843319210 $T=-19910 -20350 0 0 $X=-20820 $Y=-20780
X859 VDD 161 VDD 19 p18_CDNS_6726843319210 $T=-16780 -29620 1 0 $X=-17690 $Y=-31850
X860 VDD 160 VDD 147 p18_CDNS_6726843319210 $T=-15300 -42570 1 0 $X=-16210 $Y=-44800
X861 VDD 162 VDD 148 p18_CDNS_6726843319210 $T=-15300 -7400 0 0 $X=-16210 $Y=-7830
X862 VDD VDD 175 174 p18_CDNS_6726843319210 $T=-13400 -29620 1 0 $X=-14310 $Y=-31850
X863 VDD 181 195 145 p18_CDNS_6726843319210 $T=-10730 -33300 0 0 $X=-11640 $Y=-33730
X864 VDD 203 VDD 198 p18_CDNS_6726843319210 $T=-7840 -20350 0 0 $X=-8750 $Y=-20780
X865 VDD 230 VDD 227 p18_CDNS_6726843319210 $T=-3230 -42570 1 0 $X=-4140 $Y=-44800
X866 VDD 232 VDD 228 p18_CDNS_6726843319210 $T=-3230 -7400 0 0 $X=-4140 $Y=-7830
X867 VDD VDD 244 229 p18_CDNS_6726843319210 $T=-1290 -20350 0 0 $X=-2200 $Y=-20780
X868 VDD 252 258 226 p18_CDNS_6726843319210 $T=1340 -16670 1 0 $X=430 $Y=-18900
X869 VDD 269 VDD 260 p18_CDNS_6726843319210 $T=4230 -20350 0 0 $X=3320 $Y=-20780
X870 VDD 288 VDD 281 p18_CDNS_6726843319210 $T=8840 -42570 1 0 $X=7930 $Y=-44800
X871 VDD 290 VDD 282 p18_CDNS_6726843319210 $T=8840 -7400 0 0 $X=7930 $Y=-7830
X872 VDD 309 VDD 82 p18_CDNS_6726843319210 $T=11970 -33300 0 0 $X=11060 $Y=-33730
X873 VDD VDD 319 313 p18_CDNS_6726843319210 $T=15350 -33300 0 0 $X=14440 $Y=-33730
X874 VDD VDD 321 305 p18_CDNS_6726843319210 $T=15390 -42570 1 0 $X=14480 $Y=-44800
X875 VDD VDD 322 306 p18_CDNS_6726843319210 $T=15390 -7400 0 0 $X=14480 $Y=-7830
X876 VDD 323 VDD 316 p18_CDNS_6726843319210 $T=16300 -20350 0 0 $X=15390 $Y=-20780
X877 VDD VDD 345 338 p18_CDNS_6726843319210 $T=22810 -29620 1 0 $X=21900 $Y=-31850
X878 VDD VDD 346 331 p18_CDNS_6726843319210 $T=22850 -20350 0 0 $X=21940 $Y=-20780
X879 VDD 361 VDD 360 p18_CDNS_6726843319210 $T=28370 -20350 0 0 $X=27460 $Y=-20780
X880 VDD VDD 373 372 p18_CDNS_6726843319210 $T=34880 -29620 1 0 $X=33970 $Y=-31850
X881 VDD VDD 374 367 p18_CDNS_6726843319210 $T=34920 -20350 0 0 $X=34010 $Y=-20780
X882 VDD 377 VDD 376 p18_CDNS_6726843319210 $T=40440 -20350 0 0 $X=39530 $Y=-20780
X883 VDD VDD 383 382 p18_CDNS_6726843319210 $T=46950 -29620 1 0 $X=46040 $Y=-31850
X884 VDD VDD 384 379 p18_CDNS_6726843319210 $T=46990 -20350 0 0 $X=46080 $Y=-20780
X885 VDD 389 VDD 386 p18_CDNS_6726843319210 $T=52510 -20350 0 0 $X=51600 $Y=-20780
X886 VDD VDD 395 394 p18_CDNS_6726843319210 $T=59020 -29620 1 0 $X=58110 $Y=-31850
X887 VDD VDD 396 391 p18_CDNS_6726843319210 $T=59060 -20350 0 0 $X=58150 $Y=-20780
X888 VDD 182 196 25 146 ICV_4 $T=-12170 -16670 1 0 $X=-13080 $Y=-18900
X889 VDD 231 242 52 197 ICV_4 $T=-4710 -29620 1 0 $X=-5620 $Y=-31850
X890 VDD 251 257 63 225 ICV_4 $T=-100 -33300 0 0 $X=-1010 $Y=-33730
X891 VDD 310 314 83 280 ICV_4 $T=11970 -16670 1 0 $X=11060 $Y=-18900
X892 VDD 332 338 98 315 ICV_4 $T=19430 -29620 1 0 $X=18520 $Y=-31850
X893 VDD 368 372 117 359 ICV_4 $T=31500 -29620 1 0 $X=30590 $Y=-31850
X894 VDD 380 382 122 375 ICV_4 $T=43570 -29620 1 0 $X=42660 $Y=-31850
X895 VDD 392 394 127 385 ICV_4 $T=55640 -29620 1 0 $X=54730 $Y=-31850
X896 GND 143 12 n18_CDNS_6726843319211 $T=-18510 -26735 1 0 $X=-19210 $Y=-27305
X897 GND 145 20 n18_CDNS_6726843319211 $T=-13900 -36185 0 0 $X=-14600 $Y=-38325
X898 GND 146 21 n18_CDNS_6726843319211 $T=-13900 -13785 1 0 $X=-14600 $Y=-14355
X899 GND 197 35 n18_CDNS_6726843319211 $T=-6440 -26735 1 0 $X=-7140 $Y=-27305
X900 GND 225 55 n18_CDNS_6726843319211 $T=-1830 -36185 0 0 $X=-2530 $Y=-38325
X901 GND 226 56 n18_CDNS_6726843319211 $T=-1830 -13785 1 0 $X=-2530 $Y=-14355
X902 GND 259 68 n18_CDNS_6726843319211 $T=5630 -26735 1 0 $X=4930 $Y=-27305
X903 GND 279 80 n18_CDNS_6726843319211 $T=10240 -36185 0 0 $X=9540 $Y=-38325
X904 GND 280 81 n18_CDNS_6726843319211 $T=10240 -13785 1 0 $X=9540 $Y=-14355
X905 GND 315 95 n18_CDNS_6726843319211 $T=17700 -26735 1 0 $X=17000 $Y=-27305
X906 GND 359 114 n18_CDNS_6726843319211 $T=29770 -26735 1 0 $X=29070 $Y=-27305
X907 GND 375 121 n18_CDNS_6726843319211 $T=41840 -26735 1 0 $X=41140 $Y=-27305
X908 GND 385 126 n18_CDNS_6726843319211 $T=53910 -26735 1 0 $X=53210 $Y=-27305
X909 13 145 48 GND n18_CDNS_672684331929 $T=-18120 -36305 0 0 $X=-18780 $Y=-36655
X910 14 146 49 GND n18_CDNS_672684331929 $T=-18120 -13665 1 0 $X=-18780 $Y=-14455
X911 29 197 65 GND n18_CDNS_672684331929 $T=-10660 -26615 1 0 $X=-11320 $Y=-27405
X912 36 225 75 GND n18_CDNS_672684331929 $T=-6050 -36305 0 0 $X=-6710 $Y=-36655
X913 37 226 76 GND n18_CDNS_672684331929 $T=-6050 -13665 1 0 $X=-6710 $Y=-14455
X914 62 259 88 GND n18_CDNS_672684331929 $T=1410 -26615 1 0 $X=750 $Y=-27405
X915 71 279 285 GND n18_CDNS_672684331929 $T=6020 -36305 0 0 $X=5360 $Y=-36655
X916 72 280 286 GND n18_CDNS_672684331929 $T=6020 -13665 1 0 $X=5360 $Y=-14455
X917 85 315 109 GND n18_CDNS_672684331929 $T=13480 -26615 1 0 $X=12820 $Y=-27405
X918 106 359 120 GND n18_CDNS_672684331929 $T=25550 -26615 1 0 $X=24890 $Y=-27405
X919 119 375 125 GND n18_CDNS_672684331929 $T=37620 -26615 1 0 $X=36960 $Y=-27405
X920 124 385 388 GND n18_CDNS_672684331929 $T=49690 -26615 1 0 $X=49030 $Y=-27405
X921 GND 160 15 147 13 36 ICV_5 $T=-17830 -39565 0 180 $X=-18670 $Y=-40355
X922 GND 162 16 148 14 37 ICV_5 $T=-17830 -10405 1 180 $X=-18670 $Y=-12425
X923 GND O7 176 203 30 198 29 62 ICV_6 $T=-12420 -23355 1 180 $X=-13260 $Y=-25375
X924 GND 52 201 230 48 227 36 71 ICV_6 $T=-7810 -39565 0 180 $X=-8650 $Y=-40355
X925 GND 35 202 232 49 228 37 72 ICV_6 $T=-7810 -10405 1 180 $X=-8650 $Y=-12425
X926 GND O6 244 269 65 260 62 85 ICV_6 $T=-350 -23355 1 180 $X=-1190 $Y=-25375
X927 GND 78 267 288 75 281 71 283 ICV_6 $T=4260 -39565 0 180 $X=3420 $Y=-40355
X928 GND 68 268 290 76 282 72 284 ICV_6 $T=4260 -10405 1 180 $X=3420 $Y=-12425
X929 GND O5 298 323 88 316 85 106 ICV_6 $T=11720 -23355 1 180 $X=10880 $Y=-25375
X930 GND O4 346 361 109 360 106 119 ICV_6 $T=23790 -23355 1 180 $X=22950 $Y=-25375
X931 GND O3 374 377 120 376 119 124 ICV_6 $T=35860 -23355 1 180 $X=35020 $Y=-25375
X932 GND O2 384 389 125 386 124 387 ICV_6 $T=47930 -23355 1 180 $X=47090 $Y=-25375
X933 GND 134 133 A2 A3 8 17 B3 ICV_8 $T=-20670 -68080 1 0 $X=-21370 $Y=-68650
X934 GND 136 135 A0 A1 77 59 B3 ICV_8 $T=-20670 -61460 1 0 $X=-21370 $Y=-62030
X935 GND 138 137 Y1 Y0 60 79 X3 ICV_8 $T=-20670 9910 1 0 $X=-21370 $Y=9340
X936 GND 140 139 Y3 Y2 18 9 X3 ICV_8 $T=-20670 16530 1 0 $X=-21370 $Y=15960
X937 GND 166 165 A2 A3 57 22 B2 ICV_8 $T=-15820 -68080 1 0 $X=-16520 $Y=-68650
X938 GND 168 167 A0 A1 104 86 B2 ICV_8 $T=-15820 -61460 1 0 $X=-16520 $Y=-62030
X939 GND 170 169 Y1 Y0 87 105 X2 ICV_8 $T=-15820 9910 1 0 $X=-16520 $Y=9340
X940 GND 172 171 Y3 Y2 23 58 X2 ICV_8 $T=-15820 16530 1 0 $X=-16520 $Y=15960
X941 GND 188 187 A2 A3 53 46 B1 ICV_8 $T=-10970 -68080 1 0 $X=-11670 $Y=-68650
X942 GND 190 189 A0 A1 112 31 B1 ICV_8 $T=-10970 -61460 1 0 $X=-11670 $Y=-62030
X943 GND 192 191 Y1 Y0 32 113 X1 ICV_8 $T=-10970 9910 1 0 $X=-11670 $Y=9340
X944 GND 194 193 Y3 Y2 47 54 X1 ICV_8 $T=-10970 16530 1 0 $X=-11670 $Y=15960
X945 GND 218 217 A2 A3 101 50 B0 ICV_8 $T=-6120 -68080 1 0 $X=-6820 $Y=-68650
X946 GND 220 219 A0 A1 129 115 B0 ICV_8 $T=-6120 -61460 1 0 $X=-6820 $Y=-62030
X947 GND 222 221 Y1 Y0 116 130 X0 ICV_8 $T=-6120 9910 1 0 $X=-6820 $Y=9340
X948 GND 224 223 Y3 Y2 51 102 X0 ICV_8 $T=-6120 16530 1 0 $X=-6820 $Y=15960
X949 VDD 136 B3 p18_CDNS_672684331920 $T=-20670 -58640 0 0 $X=-21580 $Y=-59070
X950 VDD 137 X3 p18_CDNS_672684331920 $T=-20670 8670 1 0 $X=-21580 $Y=7000
X951 VDD 134 135 A2 8 A1 59 B3 ICV_9 $T=-20670 -65260 0 0 $X=-21580 $Y=-65690
X952 VDD 138 139 Y1 60 Y2 9 X3 ICV_9 $T=-20670 12730 0 0 $X=-21580 $Y=12300
X953 VDD 166 167 A2 57 A1 86 B2 ICV_9 $T=-15820 -65260 0 0 $X=-16730 $Y=-65690
X954 VDD 170 171 Y1 87 Y2 58 X2 ICV_9 $T=-15820 12730 0 0 $X=-16730 $Y=12300
X955 VDD 188 189 A2 53 A1 31 B1 ICV_9 $T=-10970 -65260 0 0 $X=-11880 $Y=-65690
X956 VDD 192 193 Y1 32 Y2 54 X1 ICV_9 $T=-10970 12730 0 0 $X=-11880 $Y=12300
X957 VDD 218 219 A2 101 A1 115 B0 ICV_9 $T=-6120 -65260 0 0 $X=-7030 $Y=-65690
X958 VDD 222 223 Y1 116 Y2 102 X0 ICV_9 $T=-6120 12730 0 0 $X=-7030 $Y=12300
X959 VDD 133 A3 17 165 22 B3 B2 ICV_11 $T=-20670 -69320 1 0 $X=-21580 $Y=-70990
X960 VDD 140 Y3 18 172 23 X3 X2 ICV_11 $T=-20670 19350 0 0 $X=-21580 $Y=18920
X961 VDD 187 A3 46 217 50 B1 B0 ICV_11 $T=-10970 -69320 1 0 $X=-11880 $Y=-70990
X962 VDD 190 A0 112 220 129 B1 B0 ICV_11 $T=-10970 -58640 0 0 $X=-11880 $Y=-59070
X963 VDD 191 Y0 113 221 130 X1 X0 ICV_11 $T=-10970 8670 1 0 $X=-11880 $Y=7000
X964 VDD 194 Y3 47 224 51 X1 X0 ICV_11 $T=-10970 19350 0 0 $X=-11880 $Y=18920
.ENDS
***************************************

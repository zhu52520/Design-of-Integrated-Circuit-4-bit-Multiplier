* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673695983861 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=3.52e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673695983860 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Buffer3 X GND VDD Y
** N=5 EP=4 IP=14 FDC=4
X0 VDD 4 X p18_CDNS_673695983861 $T=5660 -9575 0 0 $X=4750 $Y=-10005
X1 VDD Y 4 p18_CDNS_673695983861 $T=7600 -9575 0 0 $X=6690 $Y=-10005
X2 GND 4 X n18_CDNS_673695983860 $T=5660 -12195 0 0 $X=5000 $Y=-13325
X3 GND Y 4 n18_CDNS_673695983860 $T=7600 -12195 0 0 $X=6940 $Y=-13325
.ENDS
***************************************

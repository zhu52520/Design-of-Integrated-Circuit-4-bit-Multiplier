* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_672748244950 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 3 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT TSPC INVQ CLK Q RST D VDD GND
** N=14 EP=7 IP=8 FDC=15
M0 GND Q INVQ GND NM L=1.8e-07 W=4.4e-07 $X=26400 $Y=-11580 $D=0
M1 Q CLK 11 GND NM L=1.8e-07 W=4.4e-07 $X=27550 $Y=-11580 $D=0
M2 GND 5 12 GND NM L=1.8e-07 W=4.4e-07 $X=29920 $Y=-11580 $D=0
M3 5 7 GND GND NM L=1.8e-07 W=4.4e-07 $X=30640 $Y=-11580 $D=0
M4 GND RST 5 GND NM L=1.8e-07 W=4.4e-07 $X=31360 $Y=-11580 $D=0
M5 GND D 7 GND NM L=1.8e-07 W=2.2e-07 $X=33340 $Y=-11460 $D=0
M6 VDD Q INVQ VDD PM L=1.8e-07 W=8.8e-07 $X=26400 $Y=-9500 $D=4
M7 Q 4 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=27120 $Y=-9500 $D=4
M8 VDD CLK 4 VDD PM L=1.8e-07 W=8.8e-07 $X=29820 $Y=-9500 $D=4
M9 13 7 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=30540 $Y=-9500 $D=4
M10 14 RST 13 VDD PM L=1.8e-07 W=8.8e-07 $X=30970 $Y=-9500 $D=4
M11 5 CLK 14 VDD PM L=1.8e-07 W=8.8e-07 $X=31400 $Y=-9500 $D=4
M12 VDD D 7 VDD PM L=1.8e-07 W=4.4e-07 $X=33340 $Y=-9060 $D=4
X13 GND GND 4 11 n18_CDNS_672748244950 $T=27120 -11580 0 0 $X=26460 $Y=-12930
X14 GND 4 CLK 12 n18_CDNS_672748244950 $T=29490 -11580 0 0 $X=28830 $Y=-12930
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_673625162810 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673625162812 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_673625162811 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6736251628113 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673625162818 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673625162819 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 5 6 n18_CDNS_673625162818 $T=0 -1660 0 0 $X=-660 $Y=-2010
X1 3 4 5 6 n18_CDNS_673625162819 $T=0 0 0 0 $X=-660 $Y=-350
.ENDS
***************************************
.SUBCKT p18_CDNS_6736251628112 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3
** N=3 EP=3 IP=8 FDC=2
X0 1 1 2 3 p18_CDNS_6736251628112 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 3 1 2 p18_CDNS_6736251628112 $T=2020 0 0 0 $X=1070 $Y=-530
.ENDS
***************************************
.SUBCKT n18_CDNS_6736251628111 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6736251628110 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 n18_CDNS_6736251628111 $T=0 0 0 0 $X=-1520 $Y=-350
X1 3 1 2 n18_CDNS_6736251628110 $T=2020 0 0 0 $X=1360 $Y=-350
.ENDS
***************************************
.SUBCKT SRAM_Col_8bit GND BIT INVBIT SAEN OUT PCEN DATA WEN VDD ADD7 ADD6 ADD5 ADD4 ADD3 ADD2 ADD1 ADD0
** N=41 EP=17 IP=128 FDC=68
M0 GND 31 OUT GND NM L=1.8e-07 W=2.2e-07 $X=36065 $Y=-70760 $D=0
M1 GND DATA 2 GND NM L=1.8e-07 W=2.2e-07 $X=36675 $Y=-76040 $D=0
M2 22 BIT 10 GND NM L=1.8e-07 W=4.4e-07 $X=36715 $Y=-67460 $D=0
M3 22 SAEN GND GND NM L=1.8e-07 W=8.8e-07 $X=36725 $Y=-69090 $D=0
M4 40 INVBIT 22 GND NM L=1.8e-07 W=4.4e-07 $X=37435 $Y=-67460 $D=0
M5 5 2 GND GND NM L=1.8e-07 W=2.2e-07 $X=37475 $Y=-76040 $D=0
M6 GND 40 31 GND NM L=1.8e-07 W=2.2e-07 $X=38085 $Y=-70760 $D=0
M7 VDD DATA 2 VDD PM L=1.8e-07 W=4.4e-07 $X=36715 $Y=-74330 $D=4
M8 VDD 10 10 VDD PM L=1.8e-07 W=3.3e-06 $X=36715 $Y=-65050 $D=4
M9 BIT PCEN INVBIT VDD PM L=1.8e-07 W=4.4e-07 $X=36945 $Y=-11560 $D=4
M10 5 2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=37435 $Y=-74330 $D=4
M11 40 10 VDD VDD PM L=1.8e-07 W=3.3e-06 $X=37435 $Y=-65050 $D=4
X12 GND 8 BIT WEN n18_CDNS_673625162810 $T=36065 -79290 0 0 $X=35405 $Y=-79640
X13 GND INVBIT 41 WEN n18_CDNS_673625162810 $T=38085 -79290 0 0 $X=37425 $Y=-79640
X14 GND 8 GND 2 n18_CDNS_673625162812 $T=36065 -82190 0 0 $X=35405 $Y=-83320
X15 GND GND 41 5 n18_CDNS_673625162812 $T=38085 -82190 0 0 $X=37425 $Y=-83320
X16 VDD OUT 31 p18_CDNS_673625162811 $T=36245 -72410 1 180 $X=35155 $Y=-73540
X17 VDD 31 40 p18_CDNS_673625162811 $T=38265 -72410 1 180 $X=37175 $Y=-73540
X18 VDD VDD BIT PCEN p18_CDNS_6736251628113 $T=36105 -9930 0 0 $X=35195 $Y=-10360
X19 VDD INVBIT VDD PCEN p18_CDNS_6736251628113 $T=38045 -9930 0 0 $X=37135 $Y=-10360
X20 INVBIT 32 BIT 11 ADD7 GND ICV_1 $T=36555 -59520 0 90 $X=35765 $Y=-60180
X21 INVBIT 33 BIT 12 ADD6 GND ICV_1 $T=36555 -53480 0 90 $X=35765 $Y=-54140
X22 INVBIT 34 BIT 13 ADD5 GND ICV_1 $T=36555 -47440 0 90 $X=35765 $Y=-48100
X23 INVBIT 35 BIT 14 ADD4 GND ICV_1 $T=36555 -41400 0 90 $X=35765 $Y=-42060
X24 INVBIT 36 BIT 15 ADD3 GND ICV_1 $T=36555 -35360 0 90 $X=35765 $Y=-36020
X25 INVBIT 37 BIT 16 ADD2 GND ICV_1 $T=36555 -29320 0 90 $X=35765 $Y=-29980
X26 INVBIT 38 BIT 17 ADD1 GND ICV_1 $T=36555 -23280 0 90 $X=35765 $Y=-23940
X27 INVBIT 39 BIT 18 ADD0 GND ICV_1 $T=36555 -17240 0 90 $X=35765 $Y=-17900
X28 VDD 11 32 ICV_2 $T=36065 -55940 0 0 $X=35115 $Y=-56470
X29 VDD 12 33 ICV_2 $T=36065 -49900 0 0 $X=35115 $Y=-50430
X30 VDD 13 34 ICV_2 $T=36065 -43860 0 0 $X=35115 $Y=-44390
X31 VDD 14 35 ICV_2 $T=36065 -37820 0 0 $X=35115 $Y=-38350
X32 VDD 15 36 ICV_2 $T=36065 -31780 0 0 $X=35115 $Y=-32310
X33 VDD 16 37 ICV_2 $T=36065 -25740 0 0 $X=35115 $Y=-26270
X34 VDD 17 38 ICV_2 $T=36065 -19700 0 0 $X=35115 $Y=-20230
X35 VDD 18 39 ICV_2 $T=36065 -13660 0 0 $X=35115 $Y=-14190
X36 GND 11 32 ICV_3 $T=36065 -57890 0 0 $X=34545 $Y=-58240
X37 GND 12 33 ICV_3 $T=36065 -51850 0 0 $X=34545 $Y=-52200
X38 GND 13 34 ICV_3 $T=36065 -45810 0 0 $X=34545 $Y=-46160
X39 GND 14 35 ICV_3 $T=36065 -39770 0 0 $X=34545 $Y=-40120
X40 GND 15 36 ICV_3 $T=36065 -33730 0 0 $X=34545 $Y=-34080
X41 GND 16 37 ICV_3 $T=36065 -27690 0 0 $X=34545 $Y=-28040
X42 GND 17 38 ICV_3 $T=36065 -21650 0 0 $X=34545 $Y=-22000
X43 GND 18 39 ICV_3 $T=36065 -15610 0 0 $X=34545 $Y=-15960
.ENDS
***************************************

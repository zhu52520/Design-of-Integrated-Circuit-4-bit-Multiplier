* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_673633562711 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 3 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT NOR3 VDD A B GND VOUT C
** N=8 EP=6 IP=6 FDC=6
M0 VOUT B GND GND NM L=1.8e-07 W=2.2e-07 $X=-6400 $Y=530 $D=0
M1 7 A VDD VDD PM L=1.8e-07 W=1.32e-06 $X=-7200 $Y=2700 $D=4
M2 8 B 7 VDD PM L=1.8e-07 W=1.32e-06 $X=-6770 $Y=2700 $D=4
M3 VOUT C 8 VDD PM L=1.8e-07 W=1.32e-06 $X=-6340 $Y=2700 $D=4
X4 GND VOUT A n18_CDNS_673633562711 $T=-7200 530 0 0 $X=-7900 $Y=-610
X5 GND VOUT C n18_CDNS_673633562711 $T=-5600 530 0 0 $X=-6300 $Y=-610
.ENDS
***************************************

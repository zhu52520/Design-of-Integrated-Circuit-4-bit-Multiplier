* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673614678735 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT SA_v2 GND INVBIT BIT VDD SAEN OUT
** N=10 EP=6 IP=8 FDC=9
M0 5 4 GND GND NM L=1.8e-07 W=2.2e-07 $X=-9730 $Y=-2800 $D=0
M1 6 INVBIT 4 GND NM L=1.8e-07 W=4.4e-07 $X=-9080 $Y=500 $D=0
M2 6 SAEN GND GND NM L=1.8e-07 W=8.8e-07 $X=-9070 $Y=-1130 $D=0
M3 9 BIT 6 GND NM L=1.8e-07 W=4.4e-07 $X=-8360 $Y=500 $D=0
M4 OUT 5 GND GND NM L=1.8e-07 W=2.2e-07 $X=-7710 $Y=-2800 $D=0
M5 VDD 9 4 VDD PM L=1.8e-07 W=3.3e-06 $X=-9080 $Y=2910 $D=4
M6 9 9 VDD VDD PM L=1.8e-07 W=3.3e-06 $X=-8360 $Y=2910 $D=4
X7 VDD 5 4 p18_CDNS_673614678735 $T=-9730 -4450 0 0 $X=-10640 $Y=-5580
X8 VDD OUT 5 p18_CDNS_673614678735 $T=-7710 -4450 0 0 $X=-8620 $Y=-5580
.ENDS
***************************************

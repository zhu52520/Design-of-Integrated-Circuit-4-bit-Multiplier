* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_6738901947925 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947922 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 1 3 2 1 PM L=1.8e-07 W=3.3e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947929 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947921 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947923 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947918 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 5 6 n18_CDNS_6738901947923 $T=0 -1660 0 0 $X=-660 $Y=-2010
X1 3 4 5 6 n18_CDNS_6738901947918 $T=0 0 0 0 $X=-660 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947916 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947917 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=16 FDC=4
X0 1 2 1 6 n18_CDNS_6738901947916 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 1 3 7 n18_CDNS_6738901947916 $T=2020 0 0 0 $X=1360 $Y=-1130
X2 1 2 4 8 n18_CDNS_6738901947917 $T=0 2900 0 0 $X=-660 $Y=2550
X3 1 5 3 8 n18_CDNS_6738901947917 $T=2020 2900 0 0 $X=1360 $Y=2550
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=8
X0 1 2 5 3 4 10 12 11 ICV_2 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 9 7 8 13 14 11 ICV_2 $T=4460 0 0 0 $X=3800 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194795 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4
** N=5 EP=4 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_673890194795 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 1 4 p18_CDNS_673890194795 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6
** N=7 EP=6 IP=10 FDC=4
X0 1 2 3 6 ICV_4 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 6 ICV_4 $T=4460 0 0 0 $X=3550 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947920 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4
** N=5 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_6738901947920 $T=-2020 0 0 0 $X=-2930 $Y=-1130
X1 1 3 2 p18_CDNS_6738901947920 $T=0 0 0 0 $X=-910 $Y=-1130
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947924 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947919 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_6738901947924 $T=-2020 0 0 0 $X=-2720 $Y=-350
X1 1 3 2 n18_CDNS_6738901947919 $T=0 0 0 0 $X=-700 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=8
X0 1 2 3 7 ICV_6 $T=-4460 0 0 0 $X=-7390 $Y=-1130
X1 1 4 5 8 ICV_6 $T=0 0 0 0 $X=-2930 $Y=-1130
X2 6 2 3 7 ICV_7 $T=-4460 1650 0 0 $X=-7180 $Y=1300
X3 6 4 5 8 ICV_7 $T=0 1650 0 0 $X=-2720 $Y=1300
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947915 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947926 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 NM L=1.8e-07 W=8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 n18_CDNS_6738901947915 $T=0 0 0 0 $X=-1520 $Y=-350
X1 3 1 2 n18_CDNS_6738901947926 $T=2020 0 0 0 $X=1360 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_9 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 4 5 ICV_9 $T=4460 0 0 0 $X=2940 $Y=-350
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947928 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3
** N=3 EP=3 IP=8 FDC=2
X0 1 1 2 3 p18_CDNS_6738901947928 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 3 1 2 p18_CDNS_6738901947928 $T=2020 0 0 0 $X=1070 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=4
X0 1 2 3 ICV_11 $T=0 0 0 0 $X=-950 $Y=-530
X1 1 4 5 ICV_11 $T=4460 0 0 0 $X=3510 $Y=-530
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=20 FDC=16
X0 1 2 3 4 5 ICV_10 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 6 7 8 9 ICV_10 $T=8920 0 0 0 $X=7400 $Y=-350
X2 10 2 3 4 5 ICV_12 $T=0 1950 0 0 $X=-950 $Y=1420
X3 10 6 7 8 9 ICV_12 $T=8920 1950 0 0 $X=7970 $Y=1420
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=20 FDC=32
X0 1 3 4 5 6 7 8 9 10 2 ICV_13 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 11 12 13 14 15 16 17 18 2 ICV_13 $T=17840 0 0 0 $X=16320 $Y=-350
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=34 EP=34 IP=36 FDC=64
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 ICV_14 $T=0 0 0 0 $X=-1520 $Y=-350
X1 1 2 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_14 $T=35680 0 0 0 $X=34160 $Y=-350
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947913 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947914 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=3.52e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673890194799 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947911 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 n18_CDNS_6738901947911 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 3 2 n18_CDNS_6738901947911 $T=1940 0 0 0 $X=1280 $Y=-1130
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947912 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
X0 1 2 4 p18_CDNS_6738901947912 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 2 p18_CDNS_6738901947912 $T=1940 0 0 0 $X=1030 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194794 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6738901947910 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4
** N=5 EP=4 IP=7 FDC=2
X0 1 3 5 p18_CDNS_673890194794 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 2 4 5 p18_CDNS_6738901947910 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_673890194798 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=2
X0 1 2 3 5 n18_CDNS_673890194799 $T=1980 -100 0 0 $X=1320 $Y=-1230
X1 1 4 5 n18_CDNS_673890194798 $T=0 0 0 0 $X=-700 $Y=-1230
.ENDS
***************************************
.SUBCKT n18_CDNS_673890194797 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673890194796 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194790 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673890194798 $T=0 0 0 0 $X=-700 $Y=-1230
X1 1 3 5 n18_CDNS_673890194798 $T=2020 0 0 0 $X=1320 $Y=-1230
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_673890194798 $T=0 -1680 1 0 $X=-700 $Y=-2250
X1 1 3 5 n18_CDNS_673890194798 $T=0 0 0 0 $X=-700 $Y=-1230
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_21 $T=0 0 0 0 $X=-700 $Y=-2250
X1 1 4 5 8 9 ICV_21 $T=2020 0 0 0 $X=1320 $Y=-2250
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X0 1 1 2 4 p18_CDNS_673890194795 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 1 3 5 p18_CDNS_673890194795 $T=0 2360 1 0 $X=-910 $Y=790
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 2 3 6 7 ICV_23 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 8 9 ICV_23 $T=2020 0 0 0 $X=1110 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8 9
** N=9 EP=9 IP=10 FDC=4
X0 1 3 4 2 7 ICV_19 $T=4040 0 0 0 $X=3340 $Y=-1230
X1 1 5 6 8 9 ICV_20 $T=0 0 0 0 $X=-700 $Y=-1230
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7
** N=8 EP=7 IP=12 FDC=3
X0 1 1 2 5 p18_CDNS_673890194795 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 1 3 6 p18_CDNS_673890194795 $T=2020 0 0 0 $X=1110 $Y=-430
X2 1 1 4 7 p18_CDNS_673890194795 $T=4040 0 0 0 $X=3130 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 p18_CDNS_673890194790 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 p18_CDNS_673890194790 $T=0 3240 1 0 $X=-910 $Y=1230
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5
** N=5 EP=5 IP=6 FDC=2
X0 1 2 4 n18_CDNS_6738901947911 $T=0 -1480 1 0 $X=-660 $Y=-2710
X1 1 3 5 n18_CDNS_6738901947911 $T=0 0 0 0 $X=-660 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=4
X0 1 2 3 6 7 ICV_28 $T=0 0 0 0 $X=-660 $Y=-2710
X1 1 4 5 2 3 ICV_28 $T=1940 0 0 0 $X=1280 $Y=-2710
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7
** N=7 EP=7 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 7 ICV_17 $T=0 5000 1 0 $X=-910 $Y=2110
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_16 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 4 5 3 ICV_16 $T=3880 0 0 0 $X=3220 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=8
X0 1 2 3 4 5 10 ICV_31 $T=0 0 0 0 $X=-660 $Y=-1130
X1 1 6 7 8 9 5 ICV_31 $T=7760 0 0 0 $X=7100 $Y=-1130
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6
** N=7 EP=6 IP=8 FDC=4
X0 1 2 3 6 ICV_17 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 5 3 ICV_17 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4 5 6 7 8 9 10
** N=11 EP=10 IP=14 FDC=8
X0 1 2 3 4 5 10 ICV_33 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 7 8 9 5 ICV_33 $T=7760 0 0 0 $X=6850 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=14 FDC=8
X0 1 2 4 3 5 10 11 ICV_30 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 6 8 7 9 4 5 ICV_30 $T=3880 0 0 0 $X=2970 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5
** N=6 EP=5 IP=10 FDC=3
X0 1 2 3 n18_CDNS_673890194798 $T=0 0 0 0 $X=-700 $Y=-1230
X1 1 3 4 6 n18_CDNS_673890194797 $T=-2230 -100 0 0 $X=-2550 $Y=-1230
X2 1 5 6 n18_CDNS_673890194796 $T=-2660 -100 0 0 $X=-3320 $Y=-1230
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194791 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194792 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 2 3 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673890194793 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6738901947927 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT BONUS3 Q4 Q5 Q6 Q7 Q8 Q3 Q2 Q1 Q0 CLK RST SEL ADD2 ADD1 ADD0 GND MODE VDD IN0 IN1
+ IN2 IN3 IN4 IN5 IN6 IN7 IN8 IN9 IN10 IN11 IN12 IN13 IN14 IN15
** N=1567 EP=34 IP=3040 FDC=3443
M0 37 77 80 GND NM L=1.8e-07 W=4.4e-07 $X=-168335 $Y=-103525 $D=0
M1 GND 79 80 GND NM L=1.8e-07 W=4.4e-07 $X=-165675 $Y=-103525 $D=0
M2 38 81 84 GND NM L=1.8e-07 W=4.4e-07 $X=-156955 $Y=-103525 $D=0
M3 GND 83 84 GND NM L=1.8e-07 W=4.4e-07 $X=-154295 $Y=-103525 $D=0
M4 41 85 88 GND NM L=1.8e-07 W=4.4e-07 $X=-145575 $Y=-103525 $D=0
M5 GND 87 88 GND NM L=1.8e-07 W=4.4e-07 $X=-142915 $Y=-103525 $D=0
M6 42 89 92 GND NM L=1.8e-07 W=4.4e-07 $X=-134195 $Y=-103525 $D=0
M7 GND 91 92 GND NM L=1.8e-07 W=4.4e-07 $X=-131535 $Y=-103525 $D=0
M8 45 93 96 GND NM L=1.8e-07 W=4.4e-07 $X=-122815 $Y=-103525 $D=0
M9 GND 95 96 GND NM L=1.8e-07 W=4.4e-07 $X=-120155 $Y=-103525 $D=0
M10 47 97 100 GND NM L=1.8e-07 W=4.4e-07 $X=-111435 $Y=-103525 $D=0
M11 GND 99 100 GND NM L=1.8e-07 W=4.4e-07 $X=-108775 $Y=-103525 $D=0
M12 49 101 104 GND NM L=1.8e-07 W=4.4e-07 $X=-100055 $Y=-103525 $D=0
M13 GND 103 104 GND NM L=1.8e-07 W=4.4e-07 $X=-97395 $Y=-103525 $D=0
M14 52 105 108 GND NM L=1.8e-07 W=4.4e-07 $X=-88675 $Y=-103525 $D=0
M15 GND 107 108 GND NM L=1.8e-07 W=4.4e-07 $X=-86015 $Y=-103525 $D=0
M16 56 109 112 GND NM L=1.8e-07 W=4.4e-07 $X=-77295 $Y=-103525 $D=0
M17 GND 111 112 GND NM L=1.8e-07 W=4.4e-07 $X=-74635 $Y=-103525 $D=0
M18 58 113 116 GND NM L=1.8e-07 W=4.4e-07 $X=-65915 $Y=-103525 $D=0
M19 GND 115 116 GND NM L=1.8e-07 W=4.4e-07 $X=-63255 $Y=-103525 $D=0
M20 62 117 120 GND NM L=1.8e-07 W=4.4e-07 $X=-54535 $Y=-103525 $D=0
M21 GND 119 120 GND NM L=1.8e-07 W=4.4e-07 $X=-51875 $Y=-103525 $D=0
M22 66 121 124 GND NM L=1.8e-07 W=4.4e-07 $X=-43155 $Y=-103525 $D=0
M23 GND 123 124 GND NM L=1.8e-07 W=4.4e-07 $X=-40495 $Y=-103525 $D=0
M24 68 125 128 GND NM L=1.8e-07 W=4.4e-07 $X=-31775 $Y=-103525 $D=0
M25 GND 127 128 GND NM L=1.8e-07 W=4.4e-07 $X=-29115 $Y=-103525 $D=0
M26 71 129 132 GND NM L=1.8e-07 W=4.4e-07 $X=-20395 $Y=-103525 $D=0
M27 GND 131 132 GND NM L=1.8e-07 W=4.4e-07 $X=-17735 $Y=-103525 $D=0
M28 74 133 136 GND NM L=1.8e-07 W=4.4e-07 $X=-9015 $Y=-103525 $D=0
M29 GND 135 136 GND NM L=1.8e-07 W=4.4e-07 $X=-6355 $Y=-103525 $D=0
M30 76 137 141 GND NM L=1.8e-07 W=4.4e-07 $X=2365 $Y=-103525 $D=0
M31 GND 140 141 GND NM L=1.8e-07 W=4.4e-07 $X=5025 $Y=-103525 $D=0
M32 405 167 14 GND NM L=1.8e-07 W=4.4e-07 $X=17320 $Y=-12965 $D=0
M33 GND 414 144 GND NM L=1.8e-07 W=2.2e-07 $X=17400 $Y=-38765 $D=0
M34 GND 148 142 GND NM L=1.8e-07 W=2.2e-07 $X=17400 $Y=-35045 $D=0
M35 GND 149 143 GND NM L=1.8e-07 W=2.2e-07 $X=17400 $Y=13035 $D=0
M36 GND 415 145 GND NM L=1.8e-07 W=2.2e-07 $X=17400 $Y=16755 $D=0
M37 406 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=-54210 $D=0
M38 407 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=-52410 $D=0
M39 408 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=-47590 $D=0
M40 409 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=-45790 $D=0
M41 157 151 142 GND NM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-25915 $D=0
M42 404 166 14 GND NM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-9265 $D=0
M43 150 152 143 GND NM L=1.8e-07 W=4.4e-07 $X=17440 $Y=3685 $D=0
M44 410 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=23780 $D=0
M45 411 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=25580 $D=0
M46 412 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=30400 $D=0
M47 413 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=17440 $Y=32200 $D=0
M48 GND 416 405 GND NM L=1.8e-07 W=4.4e-07 $X=18040 $Y=-12965 $D=0
M49 1273 146 GND GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-38865 $D=0
M50 1274 144 GND GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-35165 $D=0
M51 148 153 157 GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-25915 $D=0
M52 149 154 150 GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=3685 $D=0
M53 1275 145 GND GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=12935 $D=0
M54 1276 147 GND GND NM L=1.8e-07 W=4.4e-07 $X=18160 $Y=16635 $D=0
M55 GND 417 404 GND NM L=1.8e-07 W=4.4e-07 $X=18240 $Y=-9265 $D=0
M56 414 160 1273 GND NM L=1.8e-07 W=4.4e-07 $X=18590 $Y=-38865 $D=0
M57 148 155 1274 GND NM L=1.8e-07 W=4.4e-07 $X=18590 $Y=-35165 $D=0
M58 149 156 1275 GND NM L=1.8e-07 W=4.4e-07 $X=18590 $Y=12935 $D=0
M59 415 161 1276 GND NM L=1.8e-07 W=4.4e-07 $X=18590 $Y=16635 $D=0
M60 416 157 GND GND NM L=1.8e-07 W=2.2e-07 $X=18800 $Y=-12865 $D=0
M61 1277 150 GND GND NM L=1.8e-07 W=4.4e-07 $X=18960 $Y=-9265 $D=0
M62 417 157 1277 GND NM L=1.8e-07 W=4.4e-07 $X=19390 $Y=-9265 $D=0
M63 155 6 11 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-54210 $D=0
M64 146 6 9 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-52410 $D=0
M65 188 6 7 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-47590 $D=0
M66 205 6 8 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-45790 $D=0
M67 207 59 65 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=23780 $D=0
M68 189 59 63 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=25580 $D=0
M69 147 59 73 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=30400 $D=0
M70 156 59 70 GND NM L=1.8e-07 W=2.2e-07 $X=19460 $Y=32200 $D=0
M71 GND 150 416 GND NM L=1.8e-07 W=2.2e-07 $X=19600 $Y=-12865 $D=0
M72 418 177 151 GND NM L=1.8e-07 W=4.4e-07 $X=19990 $Y=-22215 $D=0
M73 419 178 152 GND NM L=1.8e-07 W=4.4e-07 $X=19990 $Y=-15 $D=0
M74 420 173 151 GND NM L=1.8e-07 W=4.4e-07 $X=20100 $Y=-25915 $D=0
M75 421 174 152 GND NM L=1.8e-07 W=4.4e-07 $X=20100 $Y=3685 $D=0
M76 GND 406 155 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-54210 $D=0
M77 GND 407 146 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-52410 $D=0
M78 GND 408 188 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-47590 $D=0
M79 GND 409 205 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-45790 $D=0
M80 GND 410 207 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=23780 $D=0
M81 GND 411 189 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=25580 $D=0
M82 GND 412 147 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=30400 $D=0
M83 GND 413 156 GND NM L=1.8e-07 W=2.2e-07 $X=20260 $Y=32200 $D=0
M84 427 414 422 GND NM L=1.8e-07 W=4.4e-07 $X=20530 $Y=-38865 $D=0
M85 428 148 423 GND NM L=1.8e-07 W=4.4e-07 $X=20530 $Y=-35165 $D=0
M86 429 149 424 GND NM L=1.8e-07 W=4.4e-07 $X=20530 $Y=12935 $D=0
M87 430 415 425 GND NM L=1.8e-07 W=4.4e-07 $X=20530 $Y=16635 $D=0
M88 GND 146 427 GND NM L=1.8e-07 W=4.4e-07 $X=21250 $Y=-38865 $D=0
M89 GND 144 428 GND NM L=1.8e-07 W=4.4e-07 $X=21250 $Y=-35165 $D=0
M90 GND 145 429 GND NM L=1.8e-07 W=4.4e-07 $X=21250 $Y=12935 $D=0
M91 GND 147 430 GND NM L=1.8e-07 W=4.4e-07 $X=21250 $Y=16635 $D=0
M92 444 417 426 GND NM L=1.8e-07 W=4.4e-07 $X=21330 $Y=-9265 $D=0
M93 1278 157 445 GND NM L=1.8e-07 W=4.4e-07 $X=21580 $Y=-12965 $D=0
M94 434 177 153 GND NM L=1.8e-07 W=4.4e-07 $X=21930 $Y=-22215 $D=0
M95 435 178 154 GND NM L=1.8e-07 W=4.4e-07 $X=21930 $Y=-15 $D=0
M96 427 160 GND GND NM L=1.8e-07 W=4.4e-07 $X=21970 $Y=-38865 $D=0
M97 428 155 GND GND NM L=1.8e-07 W=4.4e-07 $X=21970 $Y=-35165 $D=0
M98 429 156 GND GND NM L=1.8e-07 W=4.4e-07 $X=21970 $Y=12935 $D=0
M99 430 161 GND GND NM L=1.8e-07 W=4.4e-07 $X=21970 $Y=16635 $D=0
M100 GND 150 1278 GND NM L=1.8e-07 W=4.4e-07 $X=22010 $Y=-12965 $D=0
M101 431 173 153 GND NM L=1.8e-07 W=4.4e-07 $X=22050 $Y=-25915 $D=0
M102 GND 150 444 GND NM L=1.8e-07 W=4.4e-07 $X=22050 $Y=-9265 $D=0
M103 433 174 154 GND NM L=1.8e-07 W=4.4e-07 $X=22050 $Y=3685 $D=0
M104 436 10 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=-54210 $D=0
M105 437 10 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=-52410 $D=0
M106 438 10 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=-47590 $D=0
M107 439 10 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=-45790 $D=0
M108 440 61 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=23780 $D=0
M109 441 61 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=25580 $D=0
M110 442 61 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=30400 $D=0
M111 443 61 GND GND NM L=1.8e-07 W=2.2e-07 $X=22290 $Y=32200 $D=0
M112 GND 418 434 GND NM L=1.8e-07 W=4.4e-07 $X=22650 $Y=-22215 $D=0
M113 GND 419 435 GND NM L=1.8e-07 W=4.4e-07 $X=22650 $Y=-15 $D=0
M114 445 416 GND GND NM L=1.8e-07 W=2.2e-07 $X=22770 $Y=-12865 $D=0
M115 444 157 GND GND NM L=1.8e-07 W=4.4e-07 $X=22770 $Y=-9265 $D=0
M116 GND 420 431 GND NM L=1.8e-07 W=4.4e-07 $X=22850 $Y=-25915 $D=0
M117 GND 421 433 GND NM L=1.8e-07 W=4.4e-07 $X=22850 $Y=3685 $D=0
M118 418 162 GND GND NM L=1.8e-07 W=2.2e-07 $X=23410 $Y=-22095 $D=0
M119 419 163 GND GND NM L=1.8e-07 W=2.2e-07 $X=23410 $Y=85 $D=0
M120 1279 158 GND GND NM L=1.8e-07 W=4.4e-07 $X=23570 $Y=-25915 $D=0
M121 1280 159 GND GND NM L=1.8e-07 W=4.4e-07 $X=23570 $Y=3685 $D=0
M122 170 422 GND GND NM L=1.8e-07 W=2.2e-07 $X=23950 $Y=-38765 $D=0
M123 158 423 GND GND NM L=1.8e-07 W=2.2e-07 $X=23950 $Y=-35045 $D=0
M124 159 424 GND GND NM L=1.8e-07 W=2.2e-07 $X=23950 $Y=13035 $D=0
M125 171 425 GND GND NM L=1.8e-07 W=2.2e-07 $X=23950 $Y=16755 $D=0
M126 420 162 1279 GND NM L=1.8e-07 W=4.4e-07 $X=24000 $Y=-25915 $D=0
M127 421 163 1280 GND NM L=1.8e-07 W=4.4e-07 $X=24000 $Y=3685 $D=0
M128 GND 158 418 GND NM L=1.8e-07 W=2.2e-07 $X=24210 $Y=-22095 $D=0
M129 GND 159 419 GND NM L=1.8e-07 W=2.2e-07 $X=24210 $Y=85 $D=0
M130 160 10 11 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-54210 $D=0
M131 186 10 9 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-52410 $D=0
M132 213 10 7 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-47590 $D=0
M133 235 10 8 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-45790 $D=0
M134 236 61 65 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=23780 $D=0
M135 214 61 63 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=25580 $D=0
M136 187 61 73 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=30400 $D=0
M137 161 61 70 GND NM L=1.8e-07 W=2.2e-07 $X=24310 $Y=32200 $D=0
M138 446 445 GND GND NM L=1.8e-07 W=4.4e-07 $X=24750 $Y=-12965 $D=0
M139 447 426 GND GND NM L=1.8e-07 W=4.4e-07 $X=24750 $Y=-9265 $D=0
M140 GND 436 160 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-54210 $D=0
M141 GND 437 186 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-52410 $D=0
M142 GND 438 213 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-47590 $D=0
M143 GND 439 235 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-45790 $D=0
M144 GND 440 236 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=23780 $D=0
M145 GND 441 214 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=25580 $D=0
M146 GND 442 187 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=30400 $D=0
M147 GND 443 161 GND NM L=1.8e-07 W=2.2e-07 $X=25110 $Y=32200 $D=0
M148 16 167 446 GND NM L=1.8e-07 W=4.4e-07 $X=25510 $Y=-12965 $D=0
M149 16 166 447 GND NM L=1.8e-07 W=4.4e-07 $X=25510 $Y=-9265 $D=0
M150 GND 486 164 GND NM L=1.8e-07 W=4.4e-07 $X=25930 $Y=-38865 $D=0
M151 GND 487 165 GND NM L=1.8e-07 W=4.4e-07 $X=25930 $Y=16635 $D=0
M152 454 420 449 GND NM L=1.8e-07 W=4.4e-07 $X=25940 $Y=-25915 $D=0
M153 455 421 450 GND NM L=1.8e-07 W=4.4e-07 $X=25940 $Y=3685 $D=0
M154 GND 456 162 GND NM L=1.8e-07 W=2.2e-07 $X=25970 $Y=-35045 $D=0
M155 GND 457 163 GND NM L=1.8e-07 W=2.2e-07 $X=25970 $Y=13035 $D=0
M156 1281 162 466 GND NM L=1.8e-07 W=4.4e-07 $X=26190 $Y=-22215 $D=0
M157 1282 163 467 GND NM L=1.8e-07 W=4.4e-07 $X=26190 $Y=-15 $D=0
M158 GND 158 1281 GND NM L=1.8e-07 W=4.4e-07 $X=26620 $Y=-22215 $D=0
M159 GND 159 1282 GND NM L=1.8e-07 W=4.4e-07 $X=26620 $Y=-15 $D=0
M160 GND 158 454 GND NM L=1.8e-07 W=4.4e-07 $X=26660 $Y=-25915 $D=0
M161 GND 159 455 GND NM L=1.8e-07 W=4.4e-07 $X=26660 $Y=3685 $D=0
M162 1283 164 GND GND NM L=1.8e-07 W=4.4e-07 $X=26730 $Y=-35165 $D=0
M163 1284 165 GND GND NM L=1.8e-07 W=4.4e-07 $X=26730 $Y=12935 $D=0
M164 458 12 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=-54210 $D=0
M165 459 12 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=-52410 $D=0
M166 460 12 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=-47590 $D=0
M167 461 12 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=-45790 $D=0
M168 462 53 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=23780 $D=0
M169 463 53 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=25580 $D=0
M170 464 53 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=30400 $D=0
M171 465 53 GND GND NM L=1.8e-07 W=2.2e-07 $X=27140 $Y=32200 $D=0
M172 456 170 1283 GND NM L=1.8e-07 W=4.4e-07 $X=27160 $Y=-35165 $D=0
M173 457 171 1284 GND NM L=1.8e-07 W=4.4e-07 $X=27160 $Y=12935 $D=0
M174 454 162 GND GND NM L=1.8e-07 W=4.4e-07 $X=27380 $Y=-25915 $D=0
M175 466 418 GND GND NM L=1.8e-07 W=2.2e-07 $X=27380 $Y=-22095 $D=0
M176 467 419 GND GND NM L=1.8e-07 W=2.2e-07 $X=27380 $Y=85 $D=0
M177 455 163 GND GND NM L=1.8e-07 W=4.4e-07 $X=27380 $Y=3685 $D=0
M178 468 193 166 GND NM L=1.8e-07 W=4.4e-07 $X=27450 $Y=-12965 $D=0
M179 469 190 166 GND NM L=1.8e-07 W=4.4e-07 $X=27560 $Y=-9265 $D=0
M180 GND 188 480 GND NM L=1.8e-07 W=4.4e-07 $X=27870 $Y=-38865 $D=0
M181 GND 189 481 GND NM L=1.8e-07 W=4.4e-07 $X=27870 $Y=16635 $D=0
M182 1285 188 GND GND NM L=1.8e-07 W=4.4e-07 $X=28590 $Y=-38865 $D=0
M183 1286 189 GND GND NM L=1.8e-07 W=4.4e-07 $X=28590 $Y=16635 $D=0
M184 486 186 1285 GND NM L=1.8e-07 W=4.4e-07 $X=29020 $Y=-38865 $D=0
M185 487 187 1286 GND NM L=1.8e-07 W=4.4e-07 $X=29020 $Y=16635 $D=0
M186 483 456 477 GND NM L=1.8e-07 W=4.4e-07 $X=29100 $Y=-35165 $D=0
M187 484 457 478 GND NM L=1.8e-07 W=4.4e-07 $X=29100 $Y=12935 $D=0
M188 175 12 11 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-54210 $D=0
M189 182 12 9 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-52410 $D=0
M190 168 12 7 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-47590 $D=0
M191 244 12 8 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-45790 $D=0
M192 245 53 65 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=23780 $D=0
M193 169 53 63 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=25580 $D=0
M194 183 53 73 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=30400 $D=0
M195 176 53 70 GND NM L=1.8e-07 W=2.2e-07 $X=29160 $Y=32200 $D=0
M196 473 449 GND GND NM L=1.8e-07 W=4.4e-07 $X=29360 $Y=-25915 $D=0
M197 471 466 GND GND NM L=1.8e-07 W=4.4e-07 $X=29360 $Y=-22215 $D=0
M198 472 467 GND GND NM L=1.8e-07 W=4.4e-07 $X=29360 $Y=-15 $D=0
M199 474 450 GND GND NM L=1.8e-07 W=4.4e-07 $X=29360 $Y=3685 $D=0
M200 476 193 167 GND NM L=1.8e-07 W=4.4e-07 $X=29390 $Y=-12965 $D=0
M201 475 190 167 GND NM L=1.8e-07 W=4.4e-07 $X=29510 $Y=-9265 $D=0
M202 480 175 486 GND NM L=1.8e-07 W=4.4e-07 $X=29740 $Y=-38865 $D=0
M203 481 176 487 GND NM L=1.8e-07 W=4.4e-07 $X=29740 $Y=16635 $D=0
M204 GND 164 483 GND NM L=1.8e-07 W=4.4e-07 $X=29820 $Y=-35165 $D=0
M205 GND 165 484 GND NM L=1.8e-07 W=4.4e-07 $X=29820 $Y=12935 $D=0
M206 GND 458 175 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-54210 $D=0
M207 GND 459 182 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-52410 $D=0
M208 GND 460 168 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-47590 $D=0
M209 GND 461 244 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-45790 $D=0
M210 GND 462 245 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=23780 $D=0
M211 GND 463 169 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=25580 $D=0
M212 GND 464 183 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=30400 $D=0
M213 GND 465 176 GND NM L=1.8e-07 W=2.2e-07 $X=29960 $Y=32200 $D=0
M214 GND 468 476 GND NM L=1.8e-07 W=4.4e-07 $X=30110 $Y=-12965 $D=0
M215 181 173 473 GND NM L=1.8e-07 W=4.4e-07 $X=30120 $Y=-25915 $D=0
M216 181 177 471 GND NM L=1.8e-07 W=4.4e-07 $X=30120 $Y=-22215 $D=0
M217 172 178 472 GND NM L=1.8e-07 W=4.4e-07 $X=30120 $Y=-15 $D=0
M218 172 174 474 GND NM L=1.8e-07 W=4.4e-07 $X=30120 $Y=3685 $D=0
M219 GND 469 475 GND NM L=1.8e-07 W=4.4e-07 $X=30310 $Y=-9265 $D=0
M220 GND 186 480 GND NM L=1.8e-07 W=4.4e-07 $X=30460 $Y=-38865 $D=0
M221 GND 187 481 GND NM L=1.8e-07 W=4.4e-07 $X=30460 $Y=16635 $D=0
M222 483 170 GND GND NM L=1.8e-07 W=4.4e-07 $X=30540 $Y=-35165 $D=0
M223 484 171 GND GND NM L=1.8e-07 W=4.4e-07 $X=30540 $Y=12935 $D=0
M224 468 181 GND GND NM L=1.8e-07 W=2.2e-07 $X=30870 $Y=-12865 $D=0
M225 1287 172 GND GND NM L=1.8e-07 W=4.4e-07 $X=31030 $Y=-9265 $D=0
M226 1288 186 GND GND NM L=1.8e-07 W=4.4e-07 $X=31180 $Y=-38865 $D=0
M227 1289 187 GND GND NM L=1.8e-07 W=4.4e-07 $X=31180 $Y=16635 $D=0
M228 469 181 1287 GND NM L=1.8e-07 W=4.4e-07 $X=31460 $Y=-9265 $D=0
M229 1290 188 1288 GND NM L=1.8e-07 W=4.4e-07 $X=31610 $Y=-38865 $D=0
M230 1291 189 1289 GND NM L=1.8e-07 W=4.4e-07 $X=31610 $Y=16635 $D=0
M231 GND 172 468 GND NM L=1.8e-07 W=2.2e-07 $X=31670 $Y=-12865 $D=0
M232 488 13 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=-54210 $D=0
M233 489 13 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=-52410 $D=0
M234 490 13 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=-47590 $D=0
M235 491 13 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=-45790 $D=0
M236 492 54 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=23780 $D=0
M237 493 54 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=25580 $D=0
M238 494 54 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=30400 $D=0
M239 495 54 GND GND NM L=1.8e-07 W=2.2e-07 $X=31990 $Y=32200 $D=0
M240 513 175 1290 GND NM L=1.8e-07 W=4.4e-07 $X=32040 $Y=-38865 $D=0
M241 514 176 1291 GND NM L=1.8e-07 W=4.4e-07 $X=32040 $Y=16635 $D=0
M242 496 203 173 GND NM L=1.8e-07 W=4.4e-07 $X=32060 $Y=-22215 $D=0
M243 497 204 174 GND NM L=1.8e-07 W=4.4e-07 $X=32060 $Y=-15 $D=0
M244 498 199 173 GND NM L=1.8e-07 W=4.4e-07 $X=32170 $Y=-25915 $D=0
M245 499 200 174 GND NM L=1.8e-07 W=4.4e-07 $X=32170 $Y=3685 $D=0
M246 184 477 GND GND NM L=1.8e-07 W=2.2e-07 $X=32520 $Y=-35045 $D=0
M247 185 478 GND GND NM L=1.8e-07 W=2.2e-07 $X=32520 $Y=13035 $D=0
M248 506 486 513 GND NM L=1.8e-07 W=4.4e-07 $X=32760 $Y=-38865 $D=0
M249 507 487 514 GND NM L=1.8e-07 W=4.4e-07 $X=32760 $Y=16635 $D=0
M250 512 469 501 GND NM L=1.8e-07 W=4.4e-07 $X=33400 $Y=-9265 $D=0
M251 GND 175 506 GND NM L=1.8e-07 W=4.4e-07 $X=33480 $Y=-38865 $D=0
M252 GND 176 507 GND NM L=1.8e-07 W=4.4e-07 $X=33480 $Y=16635 $D=0
M253 1292 181 515 GND NM L=1.8e-07 W=4.4e-07 $X=33650 $Y=-12965 $D=0
M254 509 203 177 GND NM L=1.8e-07 W=4.4e-07 $X=34000 $Y=-22215 $D=0
M255 510 204 178 GND NM L=1.8e-07 W=4.4e-07 $X=34000 $Y=-15 $D=0
M256 179 13 11 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-54210 $D=0
M257 232 13 9 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-52410 $D=0
M258 250 13 7 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-47590 $D=0
M259 278 13 8 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-45790 $D=0
M260 283 54 65 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=23780 $D=0
M261 251 54 63 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=25580 $D=0
M262 233 54 73 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=30400 $D=0
M263 180 54 70 GND NM L=1.8e-07 W=2.2e-07 $X=34010 $Y=32200 $D=0
M264 GND 172 1292 GND NM L=1.8e-07 W=4.4e-07 $X=34080 $Y=-12965 $D=0
M265 502 199 177 GND NM L=1.8e-07 W=4.4e-07 $X=34120 $Y=-25915 $D=0
M266 GND 172 512 GND NM L=1.8e-07 W=4.4e-07 $X=34120 $Y=-9265 $D=0
M267 504 200 178 GND NM L=1.8e-07 W=4.4e-07 $X=34120 $Y=3685 $D=0
M268 506 188 GND GND NM L=1.8e-07 W=4.4e-07 $X=34200 $Y=-38865 $D=0
M269 507 189 GND GND NM L=1.8e-07 W=4.4e-07 $X=34200 $Y=16635 $D=0
M270 GND 537 191 GND NM L=1.8e-07 W=4.4e-07 $X=34500 $Y=-35165 $D=0
M271 GND 538 192 GND NM L=1.8e-07 W=4.4e-07 $X=34500 $Y=12935 $D=0
M272 GND 496 509 GND NM L=1.8e-07 W=4.4e-07 $X=34720 $Y=-22215 $D=0
M273 GND 497 510 GND NM L=1.8e-07 W=4.4e-07 $X=34720 $Y=-15 $D=0
M274 GND 488 179 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-54210 $D=0
M275 GND 489 232 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-52410 $D=0
M276 GND 490 250 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-47590 $D=0
M277 GND 491 278 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-45790 $D=0
M278 GND 492 283 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=23780 $D=0
M279 GND 493 251 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=25580 $D=0
M280 GND 494 233 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=30400 $D=0
M281 GND 495 180 GND NM L=1.8e-07 W=2.2e-07 $X=34810 $Y=32200 $D=0
M282 515 468 GND GND NM L=1.8e-07 W=2.2e-07 $X=34840 $Y=-12865 $D=0
M283 512 181 GND GND NM L=1.8e-07 W=4.4e-07 $X=34840 $Y=-9265 $D=0
M284 GND 186 506 GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=-38865 $D=0
M285 GND 498 502 GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=-25915 $D=0
M286 GND 499 504 GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=3685 $D=0
M287 GND 187 507 GND NM L=1.8e-07 W=4.4e-07 $X=34920 $Y=16635 $D=0
M288 496 191 GND GND NM L=1.8e-07 W=2.2e-07 $X=35480 $Y=-22095 $D=0
M289 497 192 GND GND NM L=1.8e-07 W=2.2e-07 $X=35480 $Y=85 $D=0
M290 194 513 GND GND NM L=1.8e-07 W=4.4e-07 $X=35640 $Y=-38865 $D=0
M291 1293 184 GND GND NM L=1.8e-07 W=4.4e-07 $X=35640 $Y=-25915 $D=0
M292 1294 185 GND GND NM L=1.8e-07 W=4.4e-07 $X=35640 $Y=3685 $D=0
M293 195 514 GND GND NM L=1.8e-07 W=4.4e-07 $X=35640 $Y=16635 $D=0
M294 498 191 1293 GND NM L=1.8e-07 W=4.4e-07 $X=36070 $Y=-25915 $D=0
M295 499 192 1294 GND NM L=1.8e-07 W=4.4e-07 $X=36070 $Y=3685 $D=0
M296 GND 184 496 GND NM L=1.8e-07 W=2.2e-07 $X=36280 $Y=-22095 $D=0
M297 GND 185 497 GND NM L=1.8e-07 W=2.2e-07 $X=36280 $Y=85 $D=0
M298 GND 197 519 GND NM L=1.8e-07 W=4.4e-07 $X=36440 $Y=-35165 $D=0
M299 GND 198 522 GND NM L=1.8e-07 W=4.4e-07 $X=36440 $Y=12935 $D=0
M300 517 515 GND GND NM L=1.8e-07 W=4.4e-07 $X=36820 $Y=-12965 $D=0
M301 518 501 GND GND NM L=1.8e-07 W=4.4e-07 $X=36820 $Y=-9265 $D=0
M302 1295 197 GND GND NM L=1.8e-07 W=4.4e-07 $X=37160 $Y=-35165 $D=0
M303 1296 198 GND GND NM L=1.8e-07 W=4.4e-07 $X=37160 $Y=12935 $D=0
M304 18 193 517 GND NM L=1.8e-07 W=4.4e-07 $X=37580 $Y=-12965 $D=0
M305 18 190 518 GND NM L=1.8e-07 W=4.4e-07 $X=37580 $Y=-9265 $D=0
M306 537 201 1295 GND NM L=1.8e-07 W=4.4e-07 $X=37590 $Y=-35165 $D=0
M307 538 202 1296 GND NM L=1.8e-07 W=4.4e-07 $X=37590 $Y=12935 $D=0
M308 GND 528 201 GND NM L=1.8e-07 W=2.2e-07 $X=37620 $Y=-38765 $D=0
M309 GND 529 202 GND NM L=1.8e-07 W=2.2e-07 $X=37620 $Y=16755 $D=0
M310 530 498 524 GND NM L=1.8e-07 W=4.4e-07 $X=38010 $Y=-25915 $D=0
M311 531 499 525 GND NM L=1.8e-07 W=4.4e-07 $X=38010 $Y=3685 $D=0
M312 1297 191 532 GND NM L=1.8e-07 W=4.4e-07 $X=38260 $Y=-22215 $D=0
M313 1298 192 533 GND NM L=1.8e-07 W=4.4e-07 $X=38260 $Y=-15 $D=0
M314 519 194 537 GND NM L=1.8e-07 W=4.4e-07 $X=38310 $Y=-35165 $D=0
M315 522 195 538 GND NM L=1.8e-07 W=4.4e-07 $X=38310 $Y=12935 $D=0
M316 1299 182 GND GND NM L=1.8e-07 W=4.4e-07 $X=38380 $Y=-38865 $D=0
M317 1300 183 GND GND NM L=1.8e-07 W=4.4e-07 $X=38380 $Y=16635 $D=0
M318 GND 184 1297 GND NM L=1.8e-07 W=4.4e-07 $X=38690 $Y=-22215 $D=0
M319 GND 185 1298 GND NM L=1.8e-07 W=4.4e-07 $X=38690 $Y=-15 $D=0
M320 GND 184 530 GND NM L=1.8e-07 W=4.4e-07 $X=38730 $Y=-25915 $D=0
M321 GND 185 531 GND NM L=1.8e-07 W=4.4e-07 $X=38730 $Y=3685 $D=0
M322 528 179 1299 GND NM L=1.8e-07 W=4.4e-07 $X=38810 $Y=-38865 $D=0
M323 529 180 1300 GND NM L=1.8e-07 W=4.4e-07 $X=38810 $Y=16635 $D=0
M324 GND 201 519 GND NM L=1.8e-07 W=4.4e-07 $X=39030 $Y=-35165 $D=0
M325 GND 202 522 GND NM L=1.8e-07 W=4.4e-07 $X=39030 $Y=12935 $D=0
M326 530 191 GND GND NM L=1.8e-07 W=4.4e-07 $X=39450 $Y=-25915 $D=0
M327 532 496 GND GND NM L=1.8e-07 W=2.2e-07 $X=39450 $Y=-22095 $D=0
M328 533 497 GND GND NM L=1.8e-07 W=2.2e-07 $X=39450 $Y=85 $D=0
M329 531 192 GND GND NM L=1.8e-07 W=4.4e-07 $X=39450 $Y=3685 $D=0
M330 534 215 190 GND NM L=1.8e-07 W=4.4e-07 $X=39520 $Y=-12965 $D=0
M331 535 212 190 GND NM L=1.8e-07 W=4.4e-07 $X=39630 $Y=-9265 $D=0
M332 1301 201 GND GND NM L=1.8e-07 W=4.4e-07 $X=39750 $Y=-35165 $D=0
M333 1302 202 GND GND NM L=1.8e-07 W=4.4e-07 $X=39750 $Y=12935 $D=0
M334 1303 197 1301 GND NM L=1.8e-07 W=4.4e-07 $X=40180 $Y=-35165 $D=0
M335 1304 198 1302 GND NM L=1.8e-07 W=4.4e-07 $X=40180 $Y=12935 $D=0
M336 554 194 1303 GND NM L=1.8e-07 W=4.4e-07 $X=40610 $Y=-35165 $D=0
M337 555 195 1304 GND NM L=1.8e-07 W=4.4e-07 $X=40610 $Y=12935 $D=0
M338 547 528 539 GND NM L=1.8e-07 W=4.4e-07 $X=40750 $Y=-38865 $D=0
M339 548 529 540 GND NM L=1.8e-07 W=4.4e-07 $X=40750 $Y=16635 $D=0
M340 550 537 554 GND NM L=1.8e-07 W=4.4e-07 $X=41330 $Y=-35165 $D=0
M341 553 538 555 GND NM L=1.8e-07 W=4.4e-07 $X=41330 $Y=12935 $D=0
M342 543 524 GND GND NM L=1.8e-07 W=4.4e-07 $X=41430 $Y=-25915 $D=0
M343 541 532 GND GND NM L=1.8e-07 W=4.4e-07 $X=41430 $Y=-22215 $D=0
M344 542 533 GND GND NM L=1.8e-07 W=4.4e-07 $X=41430 $Y=-15 $D=0
M345 544 525 GND GND NM L=1.8e-07 W=4.4e-07 $X=41430 $Y=3685 $D=0
M346 546 215 193 GND NM L=1.8e-07 W=4.4e-07 $X=41460 $Y=-12965 $D=0
M347 GND 182 547 GND NM L=1.8e-07 W=4.4e-07 $X=41470 $Y=-38865 $D=0
M348 GND 183 548 GND NM L=1.8e-07 W=4.4e-07 $X=41470 $Y=16635 $D=0
M349 545 212 193 GND NM L=1.8e-07 W=4.4e-07 $X=41580 $Y=-9265 $D=0
M350 GND 194 550 GND NM L=1.8e-07 W=4.4e-07 $X=42050 $Y=-35165 $D=0
M351 GND 195 553 GND NM L=1.8e-07 W=4.4e-07 $X=42050 $Y=12935 $D=0
M352 GND 534 546 GND NM L=1.8e-07 W=4.4e-07 $X=42180 $Y=-12965 $D=0
M353 547 179 GND GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=-38865 $D=0
M354 206 199 543 GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=-25915 $D=0
M355 206 203 541 GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=-22215 $D=0
M356 196 204 542 GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=-15 $D=0
M357 196 200 544 GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=3685 $D=0
M358 548 180 GND GND NM L=1.8e-07 W=4.4e-07 $X=42190 $Y=16635 $D=0
M359 GND 535 545 GND NM L=1.8e-07 W=4.4e-07 $X=42380 $Y=-9265 $D=0
M360 550 197 GND GND NM L=1.8e-07 W=4.4e-07 $X=42770 $Y=-35165 $D=0
M361 553 198 GND GND NM L=1.8e-07 W=4.4e-07 $X=42770 $Y=12935 $D=0
M362 534 206 GND GND NM L=1.8e-07 W=2.2e-07 $X=42940 $Y=-12865 $D=0
M363 1305 196 GND GND NM L=1.8e-07 W=4.4e-07 $X=43100 $Y=-9265 $D=0
M364 GND 201 550 GND NM L=1.8e-07 W=4.4e-07 $X=43490 $Y=-35165 $D=0
M365 GND 202 553 GND NM L=1.8e-07 W=4.4e-07 $X=43490 $Y=12935 $D=0
M366 535 206 1305 GND NM L=1.8e-07 W=4.4e-07 $X=43530 $Y=-9265 $D=0
M367 GND 196 534 GND NM L=1.8e-07 W=2.2e-07 $X=43740 $Y=-12865 $D=0
M368 557 563 199 GND NM L=1.8e-07 W=4.4e-07 $X=44130 $Y=-22215 $D=0
M369 558 564 200 GND NM L=1.8e-07 W=4.4e-07 $X=44130 $Y=-15 $D=0
M370 220 539 GND GND NM L=1.8e-07 W=2.2e-07 $X=44170 $Y=-38765 $D=0
M371 221 540 GND GND NM L=1.8e-07 W=2.2e-07 $X=44170 $Y=16755 $D=0
M372 208 554 GND GND NM L=1.8e-07 W=4.4e-07 $X=44210 $Y=-35165 $D=0
M373 209 555 GND GND NM L=1.8e-07 W=4.4e-07 $X=44210 $Y=12935 $D=0
M374 559 561 199 GND NM L=1.8e-07 W=4.4e-07 $X=44240 $Y=-25915 $D=0
M375 560 562 200 GND NM L=1.8e-07 W=4.4e-07 $X=44240 $Y=3685 $D=0
M376 572 535 565 GND NM L=1.8e-07 W=4.4e-07 $X=45470 $Y=-9265 $D=0
M377 1306 206 573 GND NM L=1.8e-07 W=4.4e-07 $X=45720 $Y=-12965 $D=0
M378 570 563 203 GND NM L=1.8e-07 W=4.4e-07 $X=46070 $Y=-22215 $D=0
M379 571 564 204 GND NM L=1.8e-07 W=4.4e-07 $X=46070 $Y=-15 $D=0
M380 GND 599 210 GND NM L=1.8e-07 W=4.4e-07 $X=46150 $Y=-35165 $D=0
M381 GND 196 1306 GND NM L=1.8e-07 W=4.4e-07 $X=46150 $Y=-12965 $D=0
M382 GND 600 211 GND NM L=1.8e-07 W=4.4e-07 $X=46150 $Y=12935 $D=0
M383 GND 574 197 GND NM L=1.8e-07 W=2.2e-07 $X=46190 $Y=-38765 $D=0
M384 566 561 203 GND NM L=1.8e-07 W=4.4e-07 $X=46190 $Y=-25915 $D=0
M385 GND 196 572 GND NM L=1.8e-07 W=4.4e-07 $X=46190 $Y=-9265 $D=0
M386 568 562 204 GND NM L=1.8e-07 W=4.4e-07 $X=46190 $Y=3685 $D=0
M387 GND 575 198 GND NM L=1.8e-07 W=2.2e-07 $X=46190 $Y=16755 $D=0
M388 GND 557 570 GND NM L=1.8e-07 W=4.4e-07 $X=46790 $Y=-22215 $D=0
M389 GND 558 571 GND NM L=1.8e-07 W=4.4e-07 $X=46790 $Y=-15 $D=0
M390 573 534 GND GND NM L=1.8e-07 W=2.2e-07 $X=46910 $Y=-12865 $D=0
M391 572 206 GND GND NM L=1.8e-07 W=4.4e-07 $X=46910 $Y=-9265 $D=0
M392 1307 205 GND GND NM L=1.8e-07 W=4.4e-07 $X=46950 $Y=-38865 $D=0
M393 1308 207 GND GND NM L=1.8e-07 W=4.4e-07 $X=46950 $Y=16635 $D=0
M394 GND 559 566 GND NM L=1.8e-07 W=4.4e-07 $X=46990 $Y=-25915 $D=0
M395 GND 560 568 GND NM L=1.8e-07 W=4.4e-07 $X=46990 $Y=3685 $D=0
M396 574 213 1307 GND NM L=1.8e-07 W=4.4e-07 $X=47380 $Y=-38865 $D=0
M397 575 214 1308 GND NM L=1.8e-07 W=4.4e-07 $X=47380 $Y=16635 $D=0
M398 557 210 GND GND NM L=1.8e-07 W=2.2e-07 $X=47550 $Y=-22095 $D=0
M399 558 211 GND GND NM L=1.8e-07 W=2.2e-07 $X=47550 $Y=85 $D=0
M400 1309 208 GND GND NM L=1.8e-07 W=4.4e-07 $X=47710 $Y=-25915 $D=0
M401 1310 209 GND GND NM L=1.8e-07 W=4.4e-07 $X=47710 $Y=3685 $D=0
M402 GND 218 581 GND NM L=1.8e-07 W=4.4e-07 $X=48090 $Y=-35165 $D=0
M403 GND 219 584 GND NM L=1.8e-07 W=4.4e-07 $X=48090 $Y=12935 $D=0
M404 559 210 1309 GND NM L=1.8e-07 W=4.4e-07 $X=48140 $Y=-25915 $D=0
M405 560 211 1310 GND NM L=1.8e-07 W=4.4e-07 $X=48140 $Y=3685 $D=0
M406 GND 208 557 GND NM L=1.8e-07 W=2.2e-07 $X=48350 $Y=-22095 $D=0
M407 GND 209 558 GND NM L=1.8e-07 W=2.2e-07 $X=48350 $Y=85 $D=0
M408 1311 218 GND GND NM L=1.8e-07 W=4.4e-07 $X=48810 $Y=-35165 $D=0
M409 1312 219 GND GND NM L=1.8e-07 W=4.4e-07 $X=48810 $Y=12935 $D=0
M410 577 573 GND GND NM L=1.8e-07 W=4.4e-07 $X=48890 $Y=-12965 $D=0
M411 578 565 GND GND NM L=1.8e-07 W=4.4e-07 $X=48890 $Y=-9265 $D=0
M412 599 220 1311 GND NM L=1.8e-07 W=4.4e-07 $X=49240 $Y=-35165 $D=0
M413 600 221 1312 GND NM L=1.8e-07 W=4.4e-07 $X=49240 $Y=12935 $D=0
M414 588 574 579 GND NM L=1.8e-07 W=4.4e-07 $X=49320 $Y=-38865 $D=0
M415 589 575 580 GND NM L=1.8e-07 W=4.4e-07 $X=49320 $Y=16635 $D=0
M416 29 215 577 GND NM L=1.8e-07 W=4.4e-07 $X=49650 $Y=-12965 $D=0
M417 29 212 578 GND NM L=1.8e-07 W=4.4e-07 $X=49650 $Y=-9265 $D=0
M418 581 216 599 GND NM L=1.8e-07 W=4.4e-07 $X=49960 $Y=-35165 $D=0
M419 584 217 600 GND NM L=1.8e-07 W=4.4e-07 $X=49960 $Y=12935 $D=0
M420 GND 205 588 GND NM L=1.8e-07 W=4.4e-07 $X=50040 $Y=-38865 $D=0
M421 GND 207 589 GND NM L=1.8e-07 W=4.4e-07 $X=50040 $Y=16635 $D=0
M422 592 559 586 GND NM L=1.8e-07 W=4.4e-07 $X=50080 $Y=-25915 $D=0
M423 593 560 587 GND NM L=1.8e-07 W=4.4e-07 $X=50080 $Y=3685 $D=0
M424 1313 210 594 GND NM L=1.8e-07 W=4.4e-07 $X=50330 $Y=-22215 $D=0
M425 1314 211 595 GND NM L=1.8e-07 W=4.4e-07 $X=50330 $Y=-15 $D=0
M426 GND 220 581 GND NM L=1.8e-07 W=4.4e-07 $X=50680 $Y=-35165 $D=0
M427 GND 221 584 GND NM L=1.8e-07 W=4.4e-07 $X=50680 $Y=12935 $D=0
M428 588 213 GND GND NM L=1.8e-07 W=4.4e-07 $X=50760 $Y=-38865 $D=0
M429 GND 208 1313 GND NM L=1.8e-07 W=4.4e-07 $X=50760 $Y=-22215 $D=0
M430 GND 209 1314 GND NM L=1.8e-07 W=4.4e-07 $X=50760 $Y=-15 $D=0
M431 589 214 GND GND NM L=1.8e-07 W=4.4e-07 $X=50760 $Y=16635 $D=0
M432 GND 208 592 GND NM L=1.8e-07 W=4.4e-07 $X=50800 $Y=-25915 $D=0
M433 GND 209 593 GND NM L=1.8e-07 W=4.4e-07 $X=50800 $Y=3685 $D=0
M434 1315 220 GND GND NM L=1.8e-07 W=4.4e-07 $X=51400 $Y=-35165 $D=0
M435 1316 221 GND GND NM L=1.8e-07 W=4.4e-07 $X=51400 $Y=12935 $D=0
M436 592 210 GND GND NM L=1.8e-07 W=4.4e-07 $X=51520 $Y=-25915 $D=0
M437 594 557 GND GND NM L=1.8e-07 W=2.2e-07 $X=51520 $Y=-22095 $D=0
M438 595 558 GND GND NM L=1.8e-07 W=2.2e-07 $X=51520 $Y=85 $D=0
M439 593 211 GND GND NM L=1.8e-07 W=4.4e-07 $X=51520 $Y=3685 $D=0
M440 596 240 212 GND NM L=1.8e-07 W=4.4e-07 $X=51590 $Y=-12965 $D=0
M441 597 237 212 GND NM L=1.8e-07 W=4.4e-07 $X=51700 $Y=-9265 $D=0
M442 1317 218 1315 GND NM L=1.8e-07 W=4.4e-07 $X=51830 $Y=-35165 $D=0
M443 1318 219 1316 GND NM L=1.8e-07 W=4.4e-07 $X=51830 $Y=12935 $D=0
M444 612 216 1317 GND NM L=1.8e-07 W=4.4e-07 $X=52260 $Y=-35165 $D=0
M445 613 217 1318 GND NM L=1.8e-07 W=4.4e-07 $X=52260 $Y=12935 $D=0
M446 218 579 GND GND NM L=1.8e-07 W=2.2e-07 $X=52740 $Y=-38765 $D=0
M447 219 580 GND GND NM L=1.8e-07 W=2.2e-07 $X=52740 $Y=16755 $D=0
M448 608 599 612 GND NM L=1.8e-07 W=4.4e-07 $X=52980 $Y=-35165 $D=0
M449 611 600 613 GND NM L=1.8e-07 W=4.4e-07 $X=52980 $Y=12935 $D=0
M450 603 586 GND GND NM L=1.8e-07 W=4.4e-07 $X=53500 $Y=-25915 $D=0
M451 601 594 GND GND NM L=1.8e-07 W=4.4e-07 $X=53500 $Y=-22215 $D=0
M452 602 595 GND GND NM L=1.8e-07 W=4.4e-07 $X=53500 $Y=-15 $D=0
M453 604 587 GND GND NM L=1.8e-07 W=4.4e-07 $X=53500 $Y=3685 $D=0
M454 606 240 215 GND NM L=1.8e-07 W=4.4e-07 $X=53530 $Y=-12965 $D=0
M455 605 237 215 GND NM L=1.8e-07 W=4.4e-07 $X=53650 $Y=-9265 $D=0
M456 GND 216 608 GND NM L=1.8e-07 W=4.4e-07 $X=53700 $Y=-35165 $D=0
M457 GND 217 611 GND NM L=1.8e-07 W=4.4e-07 $X=53700 $Y=12935 $D=0
M458 GND 596 606 GND NM L=1.8e-07 W=4.4e-07 $X=54250 $Y=-12965 $D=0
M459 225 561 603 GND NM L=1.8e-07 W=4.4e-07 $X=54260 $Y=-25915 $D=0
M460 225 563 601 GND NM L=1.8e-07 W=4.4e-07 $X=54260 $Y=-22215 $D=0
M461 222 564 602 GND NM L=1.8e-07 W=4.4e-07 $X=54260 $Y=-15 $D=0
M462 222 562 604 GND NM L=1.8e-07 W=4.4e-07 $X=54260 $Y=3685 $D=0
M463 608 218 GND GND NM L=1.8e-07 W=4.4e-07 $X=54420 $Y=-35165 $D=0
M464 611 219 GND GND NM L=1.8e-07 W=4.4e-07 $X=54420 $Y=12935 $D=0
M465 GND 597 605 GND NM L=1.8e-07 W=4.4e-07 $X=54450 $Y=-9265 $D=0
M466 GND 639 216 GND NM L=1.8e-07 W=4.4e-07 $X=54720 $Y=-38865 $D=0
M467 GND 640 217 GND NM L=1.8e-07 W=4.4e-07 $X=54720 $Y=16635 $D=0
M468 596 225 GND GND NM L=1.8e-07 W=2.2e-07 $X=55010 $Y=-12865 $D=0
M469 GND 220 608 GND NM L=1.8e-07 W=4.4e-07 $X=55140 $Y=-35165 $D=0
M470 GND 221 611 GND NM L=1.8e-07 W=4.4e-07 $X=55140 $Y=12935 $D=0
M471 1319 222 GND GND NM L=1.8e-07 W=4.4e-07 $X=55170 $Y=-9265 $D=0
M472 597 225 1319 GND NM L=1.8e-07 W=4.4e-07 $X=55600 $Y=-9265 $D=0
M473 GND 222 596 GND NM L=1.8e-07 W=2.2e-07 $X=55810 $Y=-12865 $D=0
M474 229 612 GND GND NM L=1.8e-07 W=4.4e-07 $X=55860 $Y=-35165 $D=0
M475 230 613 GND GND NM L=1.8e-07 W=4.4e-07 $X=55860 $Y=12935 $D=0
M476 GND 561 563 GND NM L=1.8e-07 W=2.2e-07 $X=56240 $Y=-25815 $D=0
M477 624 20 GND GND NM L=1.8e-07 W=2.2e-07 $X=56240 $Y=-22095 $D=0
M478 625 14 GND GND NM L=1.8e-07 W=2.2e-07 $X=56240 $Y=85 $D=0
M479 GND 562 564 GND NM L=1.8e-07 W=2.2e-07 $X=56240 $Y=3805 $D=0
M480 GND 235 621 GND NM L=1.8e-07 W=4.4e-07 $X=56660 $Y=-38865 $D=0
M481 GND 236 622 GND NM L=1.8e-07 W=4.4e-07 $X=56660 $Y=16635 $D=0
M482 1320 223 GND GND NM L=1.8e-07 W=4.4e-07 $X=57000 $Y=-25915 $D=0
M483 1321 224 GND GND NM L=1.8e-07 W=4.4e-07 $X=57000 $Y=3685 $D=0
M484 1322 235 GND GND NM L=1.8e-07 W=4.4e-07 $X=57380 $Y=-38865 $D=0
M485 1323 236 GND GND NM L=1.8e-07 W=4.4e-07 $X=57380 $Y=16635 $D=0
M486 561 229 1320 GND NM L=1.8e-07 W=4.4e-07 $X=57430 $Y=-25915 $D=0
M487 562 230 1321 GND NM L=1.8e-07 W=4.4e-07 $X=57430 $Y=3685 $D=0
M488 626 597 618 GND NM L=1.8e-07 W=4.4e-07 $X=57540 $Y=-9265 $D=0
M489 1324 225 627 GND NM L=1.8e-07 W=4.4e-07 $X=57790 $Y=-12965 $D=0
M490 639 168 1322 GND NM L=1.8e-07 W=4.4e-07 $X=57810 $Y=-38865 $D=0
M491 640 169 1323 GND NM L=1.8e-07 W=4.4e-07 $X=57810 $Y=16635 $D=0
M492 GND 628 223 GND NM L=1.8e-07 W=2.2e-07 $X=57840 $Y=-35045 $D=0
M493 GND 629 224 GND NM L=1.8e-07 W=2.2e-07 $X=57840 $Y=13035 $D=0
M494 615 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=58220 $Y=-22215 $D=0
M495 GND 222 1324 GND NM L=1.8e-07 W=4.4e-07 $X=58220 $Y=-12965 $D=0
M496 616 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=58220 $Y=-15 $D=0
M497 GND 222 626 GND NM L=1.8e-07 W=4.4e-07 $X=58260 $Y=-9265 $D=0
M498 621 232 639 GND NM L=1.8e-07 W=4.4e-07 $X=58530 $Y=-38865 $D=0
M499 622 233 640 GND NM L=1.8e-07 W=4.4e-07 $X=58530 $Y=16635 $D=0
M500 1325 242 GND GND NM L=1.8e-07 W=4.4e-07 $X=58600 $Y=-35165 $D=0
M501 1326 243 GND GND NM L=1.8e-07 W=4.4e-07 $X=58600 $Y=12935 $D=0
M502 GND 624 615 GND NM L=1.8e-07 W=4.4e-07 $X=58940 $Y=-22215 $D=0
M503 GND 625 616 GND NM L=1.8e-07 W=4.4e-07 $X=58940 $Y=-15 $D=0
M504 627 596 GND GND NM L=1.8e-07 W=2.2e-07 $X=58980 $Y=-12865 $D=0
M505 626 225 GND GND NM L=1.8e-07 W=4.4e-07 $X=58980 $Y=-9265 $D=0
M506 628 238 1325 GND NM L=1.8e-07 W=4.4e-07 $X=59030 $Y=-35165 $D=0
M507 629 239 1326 GND NM L=1.8e-07 W=4.4e-07 $X=59030 $Y=12935 $D=0
M508 GND 168 621 GND NM L=1.8e-07 W=4.4e-07 $X=59250 $Y=-38865 $D=0
M509 GND 169 622 GND NM L=1.8e-07 W=4.4e-07 $X=59250 $Y=16635 $D=0
M510 635 561 631 GND NM L=1.8e-07 W=4.4e-07 $X=59370 $Y=-25915 $D=0
M511 636 562 632 GND NM L=1.8e-07 W=4.4e-07 $X=59370 $Y=3685 $D=0
M512 1327 615 GND GND NM L=1.8e-07 W=4.4e-07 $X=59660 $Y=-22215 $D=0
M513 1328 616 GND GND NM L=1.8e-07 W=4.4e-07 $X=59660 $Y=-15 $D=0
M514 1329 168 GND GND NM L=1.8e-07 W=4.4e-07 $X=59970 $Y=-38865 $D=0
M515 1330 169 GND GND NM L=1.8e-07 W=4.4e-07 $X=59970 $Y=16635 $D=0
M516 GND 223 635 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=-25915 $D=0
M517 633 CLK 1327 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=-22215 $D=0
M518 634 CLK 1328 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=-15 $D=0
M519 GND 224 636 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=3685 $D=0
M520 1331 235 1329 GND NM L=1.8e-07 W=4.4e-07 $X=60400 $Y=-38865 $D=0
M521 1332 236 1330 GND NM L=1.8e-07 W=4.4e-07 $X=60400 $Y=16635 $D=0
M522 635 229 GND GND NM L=1.8e-07 W=4.4e-07 $X=60810 $Y=-25915 $D=0
M523 636 230 GND GND NM L=1.8e-07 W=4.4e-07 $X=60810 $Y=3685 $D=0
M524 652 232 1331 GND NM L=1.8e-07 W=4.4e-07 $X=60830 $Y=-38865 $D=0
M525 653 233 1332 GND NM L=1.8e-07 W=4.4e-07 $X=60830 $Y=16635 $D=0
M526 637 627 GND GND NM L=1.8e-07 W=4.4e-07 $X=60960 $Y=-12965 $D=0
M527 638 618 GND GND NM L=1.8e-07 W=4.4e-07 $X=60960 $Y=-9265 $D=0
M528 645 628 641 GND NM L=1.8e-07 W=4.4e-07 $X=60970 $Y=-35165 $D=0
M529 646 629 642 GND NM L=1.8e-07 W=4.4e-07 $X=60970 $Y=12935 $D=0
M530 648 639 652 GND NM L=1.8e-07 W=4.4e-07 $X=61550 $Y=-38865 $D=0
M531 649 640 653 GND NM L=1.8e-07 W=4.4e-07 $X=61550 $Y=16635 $D=0
M532 GND 242 645 GND NM L=1.8e-07 W=4.4e-07 $X=61690 $Y=-35165 $D=0
M533 GND 243 646 GND NM L=1.8e-07 W=4.4e-07 $X=61690 $Y=12935 $D=0
M534 32 240 637 GND NM L=1.8e-07 W=4.4e-07 $X=61720 $Y=-12965 $D=0
M535 32 237 638 GND NM L=1.8e-07 W=4.4e-07 $X=61720 $Y=-9265 $D=0
M536 1333 CLK Q3 GND NM L=1.8e-07 W=4.4e-07 $X=62030 $Y=-22215 $D=0
M537 1334 CLK Q8 GND NM L=1.8e-07 W=4.4e-07 $X=62030 $Y=-15 $D=0
M538 GND 232 648 GND NM L=1.8e-07 W=4.4e-07 $X=62270 $Y=-38865 $D=0
M539 GND 233 649 GND NM L=1.8e-07 W=4.4e-07 $X=62270 $Y=16635 $D=0
M540 645 238 GND GND NM L=1.8e-07 W=4.4e-07 $X=62410 $Y=-35165 $D=0
M541 646 239 GND GND NM L=1.8e-07 W=4.4e-07 $X=62410 $Y=12935 $D=0
M542 GND 633 1333 GND NM L=1.8e-07 W=4.4e-07 $X=62460 $Y=-22215 $D=0
M543 GND 634 1334 GND NM L=1.8e-07 W=4.4e-07 $X=62460 $Y=-15 $D=0
M544 252 631 GND GND NM L=1.8e-07 W=2.2e-07 $X=62790 $Y=-25815 $D=0
M545 246 632 GND GND NM L=1.8e-07 W=2.2e-07 $X=62790 $Y=3805 $D=0
M546 648 235 GND GND NM L=1.8e-07 W=4.4e-07 $X=62990 $Y=-38865 $D=0
M547 649 236 GND GND NM L=1.8e-07 W=4.4e-07 $X=62990 $Y=16635 $D=0
M548 GND ADD0 234 GND NM L=1.8e-07 W=2.2e-07 $X=63050 $Y=-119495 $D=0
M549 654 260 237 GND NM L=1.8e-07 W=4.4e-07 $X=63660 $Y=-12965 $D=0
M550 GND 168 648 GND NM L=1.8e-07 W=4.4e-07 $X=63710 $Y=-38865 $D=0
M551 GND 169 649 GND NM L=1.8e-07 W=4.4e-07 $X=63710 $Y=16635 $D=0
M552 655 258 237 GND NM L=1.8e-07 W=4.4e-07 $X=63770 $Y=-9265 $D=0
M553 272 641 GND GND NM L=1.8e-07 W=2.2e-07 $X=64390 $Y=-35045 $D=0
M554 263 642 GND GND NM L=1.8e-07 W=2.2e-07 $X=64390 $Y=13035 $D=0
M555 238 652 GND GND NM L=1.8e-07 W=4.4e-07 $X=64430 $Y=-38865 $D=0
M556 239 653 GND GND NM L=1.8e-07 W=4.4e-07 $X=64430 $Y=16635 $D=0
M557 GND 241 247 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-122735 $D=0
M558 247 234 GND GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-121935 $D=0
M559 253 231 GND GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-119915 $D=0
M560 GND 241 253 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-119115 $D=0
M561 GND ADD1 254 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-115495 $D=0
M562 GND ADD1 255 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-111875 $D=0
M563 GND 241 256 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-108255 $D=0
M564 GND 241 257 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-104635 $D=0
M565 GND ADD1 248 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-101015 $D=0
M566 GND ADD1 249 GND NM L=1.8e-07 W=2.2e-07 $X=64770 $Y=-97395 $D=0
M567 664 30 GND GND NM L=1.8e-07 W=2.2e-07 $X=65160 $Y=-22095 $D=0
M568 665 16 GND GND NM L=1.8e-07 W=2.2e-07 $X=65160 $Y=85 $D=0
M569 659 260 240 GND NM L=1.8e-07 W=4.4e-07 $X=65600 $Y=-12965 $D=0
M570 658 258 240 GND NM L=1.8e-07 W=4.4e-07 $X=65720 $Y=-9265 $D=0
M571 GND 654 659 GND NM L=1.8e-07 W=4.4e-07 $X=66320 $Y=-12965 $D=0
M572 GND 666 242 GND NM L=1.8e-07 W=2.2e-07 $X=66410 $Y=-38765 $D=0
M573 GND 667 243 GND NM L=1.8e-07 W=2.2e-07 $X=66410 $Y=16755 $D=0
M574 GND 655 658 GND NM L=1.8e-07 W=4.4e-07 $X=66520 $Y=-9265 $D=0
M575 654 252 GND GND NM L=1.8e-07 W=2.2e-07 $X=67080 $Y=-12865 $D=0
M576 661 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=67140 $Y=-22215 $D=0
M577 662 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=67140 $Y=-15 $D=0
M578 1335 244 GND GND NM L=1.8e-07 W=4.4e-07 $X=67170 $Y=-38865 $D=0
M579 1336 245 GND GND NM L=1.8e-07 W=4.4e-07 $X=67170 $Y=16635 $D=0
M580 1337 246 GND GND NM L=1.8e-07 W=4.4e-07 $X=67240 $Y=-9265 $D=0
M581 666 250 1335 GND NM L=1.8e-07 W=4.4e-07 $X=67600 $Y=-38865 $D=0
M582 667 251 1336 GND NM L=1.8e-07 W=4.4e-07 $X=67600 $Y=16635 $D=0
M583 655 252 1337 GND NM L=1.8e-07 W=4.4e-07 $X=67670 $Y=-9265 $D=0
M584 GND 664 661 GND NM L=1.8e-07 W=4.4e-07 $X=67860 $Y=-22215 $D=0
M585 GND 665 662 GND NM L=1.8e-07 W=4.4e-07 $X=67860 $Y=-15 $D=0
M586 GND 246 654 GND NM L=1.8e-07 W=2.2e-07 $X=67880 $Y=-12865 $D=0
M587 1338 661 GND GND NM L=1.8e-07 W=4.4e-07 $X=68580 $Y=-22215 $D=0
M588 1339 662 GND GND NM L=1.8e-07 W=4.4e-07 $X=68580 $Y=-15 $D=0
M589 670 CLK 1338 GND NM L=1.8e-07 W=4.4e-07 $X=69010 $Y=-22215 $D=0
M590 671 CLK 1339 GND NM L=1.8e-07 W=4.4e-07 $X=69010 $Y=-15 $D=0
M591 677 666 673 GND NM L=1.8e-07 W=4.4e-07 $X=69540 $Y=-38865 $D=0
M592 678 667 674 GND NM L=1.8e-07 W=4.4e-07 $X=69540 $Y=16635 $D=0
M593 679 655 675 GND NM L=1.8e-07 W=4.4e-07 $X=69610 $Y=-9265 $D=0
M594 1340 252 680 GND NM L=1.8e-07 W=4.4e-07 $X=69860 $Y=-12965 $D=0
M595 GND 244 677 GND NM L=1.8e-07 W=4.4e-07 $X=70260 $Y=-38865 $D=0
M596 GND 245 678 GND NM L=1.8e-07 W=4.4e-07 $X=70260 $Y=16635 $D=0
M597 GND 246 1340 GND NM L=1.8e-07 W=4.4e-07 $X=70290 $Y=-12965 $D=0
M598 GND 246 679 GND NM L=1.8e-07 W=4.4e-07 $X=70330 $Y=-9265 $D=0
M599 1341 CLK Q2 GND NM L=1.8e-07 W=4.4e-07 $X=70950 $Y=-22215 $D=0
M600 1342 CLK Q7 GND NM L=1.8e-07 W=4.4e-07 $X=70950 $Y=-15 $D=0
M601 677 250 GND GND NM L=1.8e-07 W=4.4e-07 $X=70980 $Y=-38865 $D=0
M602 678 251 GND GND NM L=1.8e-07 W=4.4e-07 $X=70980 $Y=16635 $D=0
M603 680 654 GND GND NM L=1.8e-07 W=2.2e-07 $X=71050 $Y=-12865 $D=0
M604 679 252 GND GND NM L=1.8e-07 W=4.4e-07 $X=71050 $Y=-9265 $D=0
M605 GND 670 1341 GND NM L=1.8e-07 W=4.4e-07 $X=71380 $Y=-22215 $D=0
M606 GND 671 1342 GND NM L=1.8e-07 W=4.4e-07 $X=71380 $Y=-15 $D=0
M607 277 673 GND GND NM L=1.8e-07 W=2.2e-07 $X=72960 $Y=-38765 $D=0
M608 276 674 GND GND NM L=1.8e-07 W=2.2e-07 $X=72960 $Y=16755 $D=0
M609 683 680 GND GND NM L=1.8e-07 W=4.4e-07 $X=73030 $Y=-12965 $D=0
M610 684 675 GND GND NM L=1.8e-07 W=4.4e-07 $X=73030 $Y=-9265 $D=0
M611 20 260 683 GND NM L=1.8e-07 W=4.4e-07 $X=73790 $Y=-12965 $D=0
M612 20 258 684 GND NM L=1.8e-07 W=4.4e-07 $X=73790 $Y=-9265 $D=0
M613 701 34 GND GND NM L=1.8e-07 W=2.2e-07 $X=74080 $Y=-22095 $D=0
M614 702 18 GND GND NM L=1.8e-07 W=2.2e-07 $X=74080 $Y=85 $D=0
M615 699 274 258 GND NM L=1.8e-07 W=4.4e-07 $X=75730 $Y=-12965 $D=0
M616 700 273 258 GND NM L=1.8e-07 W=4.4e-07 $X=75840 $Y=-9265 $D=0
M617 695 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=76060 $Y=-22215 $D=0
M618 696 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=76060 $Y=-15 $D=0
M619 GND 701 695 GND NM L=1.8e-07 W=4.4e-07 $X=76780 $Y=-22215 $D=0
M620 GND 702 696 GND NM L=1.8e-07 W=4.4e-07 $X=76780 $Y=-15 $D=0
M621 1343 695 GND GND NM L=1.8e-07 W=4.4e-07 $X=77500 $Y=-22215 $D=0
M622 1344 696 GND GND NM L=1.8e-07 W=4.4e-07 $X=77500 $Y=-15 $D=0
M623 705 274 260 GND NM L=1.8e-07 W=4.4e-07 $X=77670 $Y=-12965 $D=0
M624 704 273 260 GND NM L=1.8e-07 W=4.4e-07 $X=77790 $Y=-9265 $D=0
M625 706 CLK 1343 GND NM L=1.8e-07 W=4.4e-07 $X=77930 $Y=-22215 $D=0
M626 707 CLK 1344 GND NM L=1.8e-07 W=4.4e-07 $X=77930 $Y=-15 $D=0
M627 715 262 GND GND NM L=1.8e-07 W=2.2e-07 $X=78350 $Y=-81965 $D=0
M628 GND 699 705 GND NM L=1.8e-07 W=4.4e-07 $X=78390 $Y=-12965 $D=0
M629 GND 700 704 GND NM L=1.8e-07 W=4.4e-07 $X=78590 $Y=-9265 $D=0
M630 699 272 GND GND NM L=1.8e-07 W=2.2e-07 $X=79150 $Y=-12865 $D=0
M631 1345 263 GND GND NM L=1.8e-07 W=4.4e-07 $X=79310 $Y=-9265 $D=0
M632 700 272 1345 GND NM L=1.8e-07 W=4.4e-07 $X=79740 $Y=-9265 $D=0
M633 1346 CLK Q1 GND NM L=1.8e-07 W=4.4e-07 $X=79870 $Y=-22215 $D=0
M634 1347 CLK Q6 GND NM L=1.8e-07 W=4.4e-07 $X=79870 $Y=-15 $D=0
M635 GND 263 699 GND NM L=1.8e-07 W=2.2e-07 $X=79950 $Y=-12865 $D=0
M636 GND 706 1346 GND NM L=1.8e-07 W=4.4e-07 $X=80300 $Y=-22215 $D=0
M637 GND 707 1347 GND NM L=1.8e-07 W=4.4e-07 $X=80300 $Y=-15 $D=0
M638 271 715 GND GND NM L=1.8e-07 W=2.2e-07 $X=80370 $Y=-81965 $D=0
M639 719 717 GND GND NM L=1.8e-07 W=8.8e-07 $X=81250 $Y=-80165 $D=0
M640 731 700 720 GND NM L=1.8e-07 W=4.4e-07 $X=81680 $Y=-9265 $D=0
M641 1348 272 732 GND NM L=1.8e-07 W=4.4e-07 $X=81930 $Y=-12965 $D=0
M642 729 271 GND GND NM L=1.8e-07 W=8.8e-07 $X=82350 $Y=-82525 $D=0
M643 GND 263 1348 GND NM L=1.8e-07 W=4.4e-07 $X=82360 $Y=-12965 $D=0
M644 GND 263 731 GND NM L=1.8e-07 W=4.4e-07 $X=82400 $Y=-9265 $D=0
M645 748 35 GND GND NM L=1.8e-07 W=2.2e-07 $X=83000 $Y=-22095 $D=0
M646 749 29 GND GND NM L=1.8e-07 W=2.2e-07 $X=83000 $Y=85 $D=0
M647 732 699 GND GND NM L=1.8e-07 W=2.2e-07 $X=83120 $Y=-12865 $D=0
M648 731 272 GND GND NM L=1.8e-07 W=4.4e-07 $X=83120 $Y=-9265 $D=0
M649 743 729 GND GND NM L=1.8e-07 W=8.8e-07 $X=84290 $Y=-82525 $D=0
M650 734 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=84980 $Y=-22215 $D=0
M651 735 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=84980 $Y=-15 $D=0
M652 745 732 GND GND NM L=1.8e-07 W=4.4e-07 $X=85100 $Y=-12965 $D=0
M653 746 720 GND GND NM L=1.8e-07 W=4.4e-07 $X=85100 $Y=-9265 $D=0
M654 GND 748 734 GND NM L=1.8e-07 W=4.4e-07 $X=85700 $Y=-22215 $D=0
M655 GND 749 735 GND NM L=1.8e-07 W=4.4e-07 $X=85700 $Y=-15 $D=0
M656 30 274 745 GND NM L=1.8e-07 W=4.4e-07 $X=85860 $Y=-12965 $D=0
M657 30 273 746 GND NM L=1.8e-07 W=4.4e-07 $X=85860 $Y=-9265 $D=0
M658 757 743 GND GND NM L=1.8e-07 W=8.8e-07 $X=86230 $Y=-82525 $D=0
M659 1349 734 GND GND NM L=1.8e-07 W=4.4e-07 $X=86420 $Y=-22215 $D=0
M660 1350 735 GND GND NM L=1.8e-07 W=4.4e-07 $X=86420 $Y=-15 $D=0
M661 760 CLK 1349 GND NM L=1.8e-07 W=4.4e-07 $X=86850 $Y=-22215 $D=0
M662 761 CLK 1350 GND NM L=1.8e-07 W=4.4e-07 $X=86850 $Y=-15 $D=0
M663 762 774 273 GND NM L=1.8e-07 W=4.4e-07 $X=87800 $Y=-12965 $D=0
M664 763 772 273 GND NM L=1.8e-07 W=4.4e-07 $X=87910 $Y=-9265 $D=0
M665 771 757 GND GND NM L=1.8e-07 W=8.8e-07 $X=88170 $Y=-82525 $D=0
M666 1351 CLK Q0 GND NM L=1.8e-07 W=4.4e-07 $X=88790 $Y=-22215 $D=0
M667 1352 CLK Q5 GND NM L=1.8e-07 W=4.4e-07 $X=88790 $Y=-15 $D=0
M668 GND 760 1351 GND NM L=1.8e-07 W=4.4e-07 $X=89220 $Y=-22215 $D=0
M669 GND 761 1352 GND NM L=1.8e-07 W=4.4e-07 $X=89220 $Y=-15 $D=0
M670 777 774 274 GND NM L=1.8e-07 W=4.4e-07 $X=89740 $Y=-12965 $D=0
M671 776 772 274 GND NM L=1.8e-07 W=4.4e-07 $X=89860 $Y=-9265 $D=0
M672 785 771 GND GND NM L=1.8e-07 W=8.8e-07 $X=90110 $Y=-82525 $D=0
M673 GND 762 777 GND NM L=1.8e-07 W=4.4e-07 $X=90460 $Y=-12965 $D=0
M674 GND 763 776 GND NM L=1.8e-07 W=4.4e-07 $X=90660 $Y=-9265 $D=0
M675 762 277 GND GND NM L=1.8e-07 W=2.2e-07 $X=91220 $Y=-12865 $D=0
M676 1353 276 GND GND NM L=1.8e-07 W=4.4e-07 $X=91380 $Y=-9265 $D=0
M677 763 277 1353 GND NM L=1.8e-07 W=4.4e-07 $X=91810 $Y=-9265 $D=0
M678 807 32 GND GND NM L=1.8e-07 W=2.2e-07 $X=91920 $Y=85 $D=0
M679 GND 276 762 GND NM L=1.8e-07 W=2.2e-07 $X=92020 $Y=-12865 $D=0
M680 797 785 GND GND NM L=1.8e-07 W=8.8e-07 $X=92050 $Y=-82525 $D=0
M681 810 763 806 GND NM L=1.8e-07 W=4.4e-07 $X=93750 $Y=-9265 $D=0
M682 789 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=93900 $Y=-15 $D=0
M683 1354 277 811 GND NM L=1.8e-07 W=4.4e-07 $X=94000 $Y=-12965 $D=0
M684 GND 276 1354 GND NM L=1.8e-07 W=4.4e-07 $X=94430 $Y=-12965 $D=0
M685 GND 276 810 GND NM L=1.8e-07 W=4.4e-07 $X=94470 $Y=-9265 $D=0
M686 GND 807 789 GND NM L=1.8e-07 W=4.4e-07 $X=94620 $Y=-15 $D=0
M687 812 788 GND GND NM L=1.8e-07 W=8.8e-07 $X=94830 $Y=-80165 $D=0
M688 811 762 GND GND NM L=1.8e-07 W=2.2e-07 $X=95190 $Y=-12865 $D=0
M689 810 277 GND GND NM L=1.8e-07 W=4.4e-07 $X=95190 $Y=-9265 $D=0
M690 1355 789 GND GND NM L=1.8e-07 W=4.4e-07 $X=95340 $Y=-15 $D=0
M691 813 CLK 1355 GND NM L=1.8e-07 W=4.4e-07 $X=95770 $Y=-15 $D=0
M692 824 271 1356 GND NM L=1.8e-07 W=4.4e-07 $X=96440 $Y=-82085 $D=0
M693 815 811 GND GND NM L=1.8e-07 W=4.4e-07 $X=97170 $Y=-12965 $D=0
M694 816 806 GND GND NM L=1.8e-07 W=4.4e-07 $X=97170 $Y=-9265 $D=0
M695 1357 CLK Q4 GND NM L=1.8e-07 W=4.4e-07 $X=97710 $Y=-15 $D=0
M696 34 774 815 GND NM L=1.8e-07 W=4.4e-07 $X=97930 $Y=-12965 $D=0
M697 34 772 816 GND NM L=1.8e-07 W=4.4e-07 $X=97930 $Y=-9265 $D=0
M698 GND 813 1357 GND NM L=1.8e-07 W=4.4e-07 $X=98140 $Y=-15 $D=0
M699 1358 CLK GND GND NM L=1.8e-07 W=4.4e-07 $X=98790 $Y=-80165 $D=0
M700 836 826 1358 GND NM L=1.8e-07 W=4.4e-07 $X=99220 $Y=-80165 $D=0
M701 GND 772 774 GND NM L=1.8e-07 W=2.2e-07 $X=99910 $Y=-9145 $D=0
M702 1359 278 GND GND NM L=1.8e-07 W=4.4e-07 $X=100670 $Y=-9265 $D=0
M703 838 828 1360 GND NM L=1.8e-07 W=4.4e-07 $X=101080 $Y=-141125 $D=0
M704 845 835 1361 GND NM L=1.8e-07 W=4.4e-07 $X=101080 $Y=-82085 $D=0
M705 772 283 1359 GND NM L=1.8e-07 W=4.4e-07 $X=101100 $Y=-9265 $D=0
M706 847 772 846 GND NM L=1.8e-07 W=4.4e-07 $X=103040 $Y=-9265 $D=0
M707 848 838 GND GND NM L=1.8e-07 W=2.2e-07 $X=103310 $Y=-141025 $D=0
M708 855 845 GND GND NM L=1.8e-07 W=2.2e-07 $X=103310 $Y=-81965 $D=0
M709 GND 278 847 GND NM L=1.8e-07 W=4.4e-07 $X=103760 $Y=-9265 $D=0
M710 847 283 GND GND NM L=1.8e-07 W=4.4e-07 $X=104480 $Y=-9265 $D=0
M711 284 848 GND GND NM L=1.8e-07 W=2.2e-07 $X=105330 $Y=-141025 $D=0
M712 291 855 GND GND NM L=1.8e-07 W=2.2e-07 $X=105330 $Y=-81965 $D=0
M713 35 846 GND GND NM L=1.8e-07 W=2.2e-07 $X=106460 $Y=-9145 $D=0
M714 294 19 GND GND NM L=1.8e-07 W=2.2e-07 $X=107350 $Y=-141025 $D=0
M715 303 MODE 262 GND NM L=1.8e-07 W=4.4e-07 $X=107470 $Y=-80165 $D=0
M716 261 279 302 GND NM L=1.8e-07 W=4.4e-07 $X=108190 $Y=-143045 $D=0
M717 262 280 303 GND NM L=1.8e-07 W=4.4e-07 $X=108190 $Y=-80165 $D=0
M718 302 281 GND GND NM L=1.8e-07 W=4.4e-07 $X=110130 $Y=-143045 $D=0
M719 303 282 GND GND NM L=1.8e-07 W=4.4e-07 $X=110130 $Y=-80165 $D=0
M720 GND 292 302 GND NM L=1.8e-07 W=4.4e-07 $X=110850 $Y=-143045 $D=0
M721 GND 293 303 GND NM L=1.8e-07 W=4.4e-07 $X=110850 $Y=-80165 $D=0
M722 866 284 313 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-141125 $D=0
M723 867 285 314 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-127805 $D=0
M724 868 286 315 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-125885 $D=0
M725 863 287 316 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-112565 $D=0
M726 864 288 317 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-110645 $D=0
M727 869 289 318 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-97325 $D=0
M728 870 290 319 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-95405 $D=0
M729 871 291 320 GND NM L=1.8e-07 W=4.4e-07 $X=112070 $Y=-82085 $D=0
M730 320 301 GND GND NM L=1.8e-07 W=4.4e-07 $X=114010 $Y=-82085 $D=0
M731 865 861 GND GND NM L=1.8e-07 W=8.8e-07 $X=114730 $Y=-143485 $D=0
M732 GND 305 313 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-141125 $D=0
M733 GND 306 314 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-127805 $D=0
M734 GND 307 315 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-125885 $D=0
M735 GND 308 316 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-112565 $D=0
M736 GND 309 317 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-110645 $D=0
M737 GND 310 318 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-97325 $D=0
M738 GND 311 319 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-95405 $D=0
M739 GND 312 320 GND NM L=1.8e-07 W=4.4e-07 $X=114730 $Y=-82085 $D=0
M740 1362 894 GND GND NM L=1.8e-07 W=4.4e-07 $X=118450 $Y=-164780 $D=0
M741 1363 895 GND GND NM L=1.8e-07 W=4.4e-07 $X=118450 $Y=-161080 $D=0
M742 7 323 1362 GND NM L=1.8e-07 W=4.4e-07 $X=118880 $Y=-164780 $D=0
M743 8 323 1363 GND NM L=1.8e-07 W=4.4e-07 $X=118880 $Y=-161080 $D=0
M744 GND 37 322 GND NM L=1.8e-07 W=2.2e-07 $X=119060 $Y=-148195 $D=0
M745 883 324 874 GND NM L=1.8e-07 W=4.4e-07 $X=119100 $Y=-139615 $D=0
M746 326 322 GND GND NM L=1.8e-07 W=2.2e-07 $X=119860 $Y=-148195 $D=0
M747 1364 323 894 GND NM L=1.8e-07 W=4.4e-07 $X=120820 $Y=-164780 $D=0
M748 1365 323 895 GND NM L=1.8e-07 W=4.4e-07 $X=120820 $Y=-161080 $D=0
M749 GND 898 1364 GND NM L=1.8e-07 W=4.4e-07 $X=121250 $Y=-164780 $D=0
M750 GND 899 1365 GND NM L=1.8e-07 W=4.4e-07 $X=121250 $Y=-161080 $D=0
M751 898 910 GND GND NM L=1.8e-07 W=4.4e-07 $X=121970 $Y=-164780 $D=0
M752 899 911 GND GND NM L=1.8e-07 W=4.4e-07 $X=121970 $Y=-161080 $D=0
M753 GND RST 898 GND NM L=1.8e-07 W=4.4e-07 $X=122690 $Y=-164780 $D=0
M754 GND RST 899 GND NM L=1.8e-07 W=4.4e-07 $X=122690 $Y=-161080 $D=0
M755 GND 38 327 GND NM L=1.8e-07 W=2.2e-07 $X=123520 $Y=-148195 $D=0
M756 909 328 900 GND NM L=1.8e-07 W=4.4e-07 $X=123560 $Y=-139615 $D=0
M757 330 327 GND GND NM L=1.8e-07 W=2.2e-07 $X=124320 $Y=-148195 $D=0
M758 GND 39 910 GND NM L=1.8e-07 W=2.2e-07 $X=124670 $Y=-164680 $D=0
M759 GND 36 911 GND NM L=1.8e-07 W=2.2e-07 $X=124670 $Y=-160960 $D=0
M760 1366 934 GND GND NM L=1.8e-07 W=4.4e-07 $X=126650 $Y=-164780 $D=0
M761 1367 935 GND GND NM L=1.8e-07 W=4.4e-07 $X=126650 $Y=-161080 $D=0
M762 11 323 1366 GND NM L=1.8e-07 W=4.4e-07 $X=127080 $Y=-164780 $D=0
M763 9 323 1367 GND NM L=1.8e-07 W=4.4e-07 $X=127080 $Y=-161080 $D=0
M764 GND 41 331 GND NM L=1.8e-07 W=2.2e-07 $X=127980 $Y=-148195 $D=0
M765 933 332 924 GND NM L=1.8e-07 W=4.4e-07 $X=128020 $Y=-139615 $D=0
M766 334 331 GND GND NM L=1.8e-07 W=2.2e-07 $X=128780 $Y=-148195 $D=0
M767 1368 323 934 GND NM L=1.8e-07 W=4.4e-07 $X=129020 $Y=-164780 $D=0
M768 1369 323 935 GND NM L=1.8e-07 W=4.4e-07 $X=129020 $Y=-161080 $D=0
M769 GND 948 1368 GND NM L=1.8e-07 W=4.4e-07 $X=129450 $Y=-164780 $D=0
M770 GND 949 1369 GND NM L=1.8e-07 W=4.4e-07 $X=129450 $Y=-161080 $D=0
M771 948 959 GND GND NM L=1.8e-07 W=4.4e-07 $X=130170 $Y=-164780 $D=0
M772 949 960 GND GND NM L=1.8e-07 W=4.4e-07 $X=130170 $Y=-161080 $D=0
M773 GND RST 948 GND NM L=1.8e-07 W=4.4e-07 $X=130890 $Y=-164780 $D=0
M774 GND RST 949 GND NM L=1.8e-07 W=4.4e-07 $X=130890 $Y=-161080 $D=0
M775 GND 42 335 GND NM L=1.8e-07 W=2.2e-07 $X=132440 $Y=-148195 $D=0
M776 961 336 950 GND NM L=1.8e-07 W=4.4e-07 $X=132480 $Y=-139615 $D=0
M777 GND 43 959 GND NM L=1.8e-07 W=2.2e-07 $X=132870 $Y=-164680 $D=0
M778 GND 40 960 GND NM L=1.8e-07 W=2.2e-07 $X=132870 $Y=-160960 $D=0
M779 338 335 GND GND NM L=1.8e-07 W=2.2e-07 $X=133240 $Y=-148195 $D=0
M780 1370 983 GND GND NM L=1.8e-07 W=4.4e-07 $X=134850 $Y=-164780 $D=0
M781 1371 984 GND GND NM L=1.8e-07 W=4.4e-07 $X=134850 $Y=-161080 $D=0
M782 12 323 1370 GND NM L=1.8e-07 W=4.4e-07 $X=135280 $Y=-164780 $D=0
M783 13 323 1371 GND NM L=1.8e-07 W=4.4e-07 $X=135280 $Y=-161080 $D=0
M784 GND 45 339 GND NM L=1.8e-07 W=2.2e-07 $X=136900 $Y=-148195 $D=0
M785 985 340 974 GND NM L=1.8e-07 W=4.4e-07 $X=136940 $Y=-139615 $D=0
M786 1372 323 983 GND NM L=1.8e-07 W=4.4e-07 $X=137220 $Y=-164780 $D=0
M787 1373 323 984 GND NM L=1.8e-07 W=4.4e-07 $X=137220 $Y=-161080 $D=0
M788 GND 997 1372 GND NM L=1.8e-07 W=4.4e-07 $X=137650 $Y=-164780 $D=0
M789 GND 998 1373 GND NM L=1.8e-07 W=4.4e-07 $X=137650 $Y=-161080 $D=0
M790 342 339 GND GND NM L=1.8e-07 W=2.2e-07 $X=137700 $Y=-148195 $D=0
M791 997 1000 GND GND NM L=1.8e-07 W=4.4e-07 $X=138370 $Y=-164780 $D=0
M792 998 1001 GND GND NM L=1.8e-07 W=4.4e-07 $X=138370 $Y=-161080 $D=0
M793 GND RST 997 GND NM L=1.8e-07 W=4.4e-07 $X=139090 $Y=-164780 $D=0
M794 GND RST 998 GND NM L=1.8e-07 W=4.4e-07 $X=139090 $Y=-161080 $D=0
M795 GND 46 1000 GND NM L=1.8e-07 W=2.2e-07 $X=141070 $Y=-164680 $D=0
M796 GND 44 1001 GND NM L=1.8e-07 W=2.2e-07 $X=141070 $Y=-160960 $D=0
M797 GND 47 343 GND NM L=1.8e-07 W=2.2e-07 $X=141360 $Y=-148195 $D=0
M798 1011 344 1002 GND NM L=1.8e-07 W=4.4e-07 $X=141400 $Y=-139615 $D=0
M799 346 343 GND GND NM L=1.8e-07 W=2.2e-07 $X=142160 $Y=-148195 $D=0
M800 1374 1024 GND GND NM L=1.8e-07 W=4.4e-07 $X=143050 $Y=-164780 $D=0
M801 1375 1025 GND GND NM L=1.8e-07 W=4.4e-07 $X=143050 $Y=-161080 $D=0
M802 6 323 1374 GND NM L=1.8e-07 W=4.4e-07 $X=143480 $Y=-164780 $D=0
M803 10 323 1375 GND NM L=1.8e-07 W=4.4e-07 $X=143480 $Y=-161080 $D=0
M804 1376 323 1024 GND NM L=1.8e-07 W=4.4e-07 $X=145420 $Y=-164780 $D=0
M805 1377 323 1025 GND NM L=1.8e-07 W=4.4e-07 $X=145420 $Y=-161080 $D=0
M806 GND 49 347 GND NM L=1.8e-07 W=2.2e-07 $X=145820 $Y=-148195 $D=0
M807 GND 1047 1376 GND NM L=1.8e-07 W=4.4e-07 $X=145850 $Y=-164780 $D=0
M808 GND 1048 1377 GND NM L=1.8e-07 W=4.4e-07 $X=145850 $Y=-161080 $D=0
M809 1035 348 1026 GND NM L=1.8e-07 W=4.4e-07 $X=145860 $Y=-139615 $D=0
M810 1047 1049 GND GND NM L=1.8e-07 W=4.4e-07 $X=146570 $Y=-164780 $D=0
M811 1048 1050 GND GND NM L=1.8e-07 W=4.4e-07 $X=146570 $Y=-161080 $D=0
M812 350 347 GND GND NM L=1.8e-07 W=2.2e-07 $X=146620 $Y=-148195 $D=0
M813 GND RST 1047 GND NM L=1.8e-07 W=4.4e-07 $X=147290 $Y=-164780 $D=0
M814 GND RST 1048 GND NM L=1.8e-07 W=4.4e-07 $X=147290 $Y=-161080 $D=0
M815 GND 51 1049 GND NM L=1.8e-07 W=2.2e-07 $X=149270 $Y=-164680 $D=0
M816 GND 48 1050 GND NM L=1.8e-07 W=2.2e-07 $X=149270 $Y=-160960 $D=0
M817 GND 52 351 GND NM L=1.8e-07 W=2.2e-07 $X=150280 $Y=-148195 $D=0
M818 1061 352 1052 GND NM L=1.8e-07 W=4.4e-07 $X=150320 $Y=-139615 $D=0
M819 354 351 GND GND NM L=1.8e-07 W=2.2e-07 $X=151080 $Y=-148195 $D=0
M820 1378 1073 GND GND NM L=1.8e-07 W=4.4e-07 $X=151250 $Y=-164780 $D=0
M821 1379 1074 GND GND NM L=1.8e-07 W=4.4e-07 $X=151250 $Y=-161080 $D=0
M822 53 323 1378 GND NM L=1.8e-07 W=4.4e-07 $X=151680 $Y=-164780 $D=0
M823 54 323 1379 GND NM L=1.8e-07 W=4.4e-07 $X=151680 $Y=-161080 $D=0
M824 1380 323 1073 GND NM L=1.8e-07 W=4.4e-07 $X=153620 $Y=-164780 $D=0
M825 1381 323 1074 GND NM L=1.8e-07 W=4.4e-07 $X=153620 $Y=-161080 $D=0
M826 GND 1095 1380 GND NM L=1.8e-07 W=4.4e-07 $X=154050 $Y=-164780 $D=0
M827 GND 1096 1381 GND NM L=1.8e-07 W=4.4e-07 $X=154050 $Y=-161080 $D=0
M828 GND 56 355 GND NM L=1.8e-07 W=2.2e-07 $X=154740 $Y=-148195 $D=0
M829 1095 1099 GND GND NM L=1.8e-07 W=4.4e-07 $X=154770 $Y=-164780 $D=0
M830 1096 1100 GND GND NM L=1.8e-07 W=4.4e-07 $X=154770 $Y=-161080 $D=0
M831 1085 356 1076 GND NM L=1.8e-07 W=4.4e-07 $X=154780 $Y=-139615 $D=0
M832 GND RST 1095 GND NM L=1.8e-07 W=4.4e-07 $X=155490 $Y=-164780 $D=0
M833 GND RST 1096 GND NM L=1.8e-07 W=4.4e-07 $X=155490 $Y=-161080 $D=0
M834 358 355 GND GND NM L=1.8e-07 W=2.2e-07 $X=155540 $Y=-148195 $D=0
M835 GND 57 1099 GND NM L=1.8e-07 W=2.2e-07 $X=157470 $Y=-164680 $D=0
M836 GND 55 1100 GND NM L=1.8e-07 W=2.2e-07 $X=157470 $Y=-160960 $D=0
M837 GND 58 359 GND NM L=1.8e-07 W=2.2e-07 $X=159200 $Y=-148195 $D=0
M838 1111 360 1102 GND NM L=1.8e-07 W=4.4e-07 $X=159240 $Y=-139615 $D=0
M839 1382 1123 GND GND NM L=1.8e-07 W=4.4e-07 $X=159450 $Y=-164780 $D=0
M840 1383 1124 GND GND NM L=1.8e-07 W=4.4e-07 $X=159450 $Y=-161080 $D=0
M841 59 323 1382 GND NM L=1.8e-07 W=4.4e-07 $X=159880 $Y=-164780 $D=0
M842 61 323 1383 GND NM L=1.8e-07 W=4.4e-07 $X=159880 $Y=-161080 $D=0
M843 362 359 GND GND NM L=1.8e-07 W=2.2e-07 $X=160000 $Y=-148195 $D=0
M844 1384 323 1123 GND NM L=1.8e-07 W=4.4e-07 $X=161820 $Y=-164780 $D=0
M845 1385 323 1124 GND NM L=1.8e-07 W=4.4e-07 $X=161820 $Y=-161080 $D=0
M846 GND 1136 1384 GND NM L=1.8e-07 W=4.4e-07 $X=162250 $Y=-164780 $D=0
M847 GND 1137 1385 GND NM L=1.8e-07 W=4.4e-07 $X=162250 $Y=-161080 $D=0
M848 1136 1148 GND GND NM L=1.8e-07 W=4.4e-07 $X=162970 $Y=-164780 $D=0
M849 1137 1149 GND GND NM L=1.8e-07 W=4.4e-07 $X=162970 $Y=-161080 $D=0
M850 GND 62 363 GND NM L=1.8e-07 W=2.2e-07 $X=163660 $Y=-148195 $D=0
M851 GND RST 1136 GND NM L=1.8e-07 W=4.4e-07 $X=163690 $Y=-164780 $D=0
M852 GND RST 1137 GND NM L=1.8e-07 W=4.4e-07 $X=163690 $Y=-161080 $D=0
M853 1135 364 1126 GND NM L=1.8e-07 W=4.4e-07 $X=163700 $Y=-139615 $D=0
M854 366 363 GND GND NM L=1.8e-07 W=2.2e-07 $X=164460 $Y=-148195 $D=0
M855 GND 64 1148 GND NM L=1.8e-07 W=2.2e-07 $X=165670 $Y=-164680 $D=0
M856 GND 60 1149 GND NM L=1.8e-07 W=2.2e-07 $X=165670 $Y=-160960 $D=0
M857 1386 1173 GND GND NM L=1.8e-07 W=4.4e-07 $X=167650 $Y=-164780 $D=0
M858 1387 1174 GND GND NM L=1.8e-07 W=4.4e-07 $X=167650 $Y=-161080 $D=0
M859 63 323 1386 GND NM L=1.8e-07 W=4.4e-07 $X=168080 $Y=-164780 $D=0
M860 65 323 1387 GND NM L=1.8e-07 W=4.4e-07 $X=168080 $Y=-161080 $D=0
M861 GND 66 367 GND NM L=1.8e-07 W=2.2e-07 $X=168120 $Y=-148195 $D=0
M862 1161 368 1152 GND NM L=1.8e-07 W=4.4e-07 $X=168160 $Y=-139615 $D=0
M863 370 367 GND GND NM L=1.8e-07 W=2.2e-07 $X=168920 $Y=-148195 $D=0
M864 1388 323 1173 GND NM L=1.8e-07 W=4.4e-07 $X=170020 $Y=-164780 $D=0
M865 1389 323 1174 GND NM L=1.8e-07 W=4.4e-07 $X=170020 $Y=-161080 $D=0
M866 GND 1177 1388 GND NM L=1.8e-07 W=4.4e-07 $X=170450 $Y=-164780 $D=0
M867 GND 1178 1389 GND NM L=1.8e-07 W=4.4e-07 $X=170450 $Y=-161080 $D=0
M868 1177 1188 GND GND NM L=1.8e-07 W=4.4e-07 $X=171170 $Y=-164780 $D=0
M869 1178 1189 GND GND NM L=1.8e-07 W=4.4e-07 $X=171170 $Y=-161080 $D=0
M870 GND RST 1177 GND NM L=1.8e-07 W=4.4e-07 $X=171890 $Y=-164780 $D=0
M871 GND RST 1178 GND NM L=1.8e-07 W=4.4e-07 $X=171890 $Y=-161080 $D=0
M872 GND 68 371 GND NM L=1.8e-07 W=2.2e-07 $X=172580 $Y=-148195 $D=0
M873 1187 372 1176 GND NM L=1.8e-07 W=4.4e-07 $X=172620 $Y=-139615 $D=0
M874 374 371 GND GND NM L=1.8e-07 W=2.2e-07 $X=173380 $Y=-148195 $D=0
M875 GND 69 1188 GND NM L=1.8e-07 W=2.2e-07 $X=173870 $Y=-164680 $D=0
M876 GND 67 1189 GND NM L=1.8e-07 W=2.2e-07 $X=173870 $Y=-160960 $D=0
M877 1390 1221 GND GND NM L=1.8e-07 W=4.4e-07 $X=175850 $Y=-164780 $D=0
M878 1391 1222 GND GND NM L=1.8e-07 W=4.4e-07 $X=175850 $Y=-161080 $D=0
M879 70 323 1390 GND NM L=1.8e-07 W=4.4e-07 $X=176280 $Y=-164780 $D=0
M880 73 323 1391 GND NM L=1.8e-07 W=4.4e-07 $X=176280 $Y=-161080 $D=0
M881 GND 71 375 GND NM L=1.8e-07 W=2.2e-07 $X=177040 $Y=-148195 $D=0
M882 1211 376 1202 GND NM L=1.8e-07 W=4.4e-07 $X=177080 $Y=-139615 $D=0
M883 378 375 GND GND NM L=1.8e-07 W=2.2e-07 $X=177840 $Y=-148195 $D=0
M884 1392 323 1221 GND NM L=1.8e-07 W=4.4e-07 $X=178220 $Y=-164780 $D=0
M885 1393 323 1222 GND NM L=1.8e-07 W=4.4e-07 $X=178220 $Y=-161080 $D=0
M886 GND 1226 1392 GND NM L=1.8e-07 W=4.4e-07 $X=178650 $Y=-164780 $D=0
M887 GND 1227 1393 GND NM L=1.8e-07 W=4.4e-07 $X=178650 $Y=-161080 $D=0
M888 1226 1237 GND GND NM L=1.8e-07 W=4.4e-07 $X=179370 $Y=-164780 $D=0
M889 1227 1238 GND GND NM L=1.8e-07 W=4.4e-07 $X=179370 $Y=-161080 $D=0
M890 GND RST 1226 GND NM L=1.8e-07 W=4.4e-07 $X=180090 $Y=-164780 $D=0
M891 GND RST 1227 GND NM L=1.8e-07 W=4.4e-07 $X=180090 $Y=-161080 $D=0
M892 GND 74 379 GND NM L=1.8e-07 W=2.2e-07 $X=181500 $Y=-148195 $D=0
M893 1239 380 1228 GND NM L=1.8e-07 W=4.4e-07 $X=181540 $Y=-139615 $D=0
M894 GND 75 1237 GND NM L=1.8e-07 W=2.2e-07 $X=182070 $Y=-164680 $D=0
M895 GND 72 1238 GND NM L=1.8e-07 W=2.2e-07 $X=182070 $Y=-160960 $D=0
M896 382 379 GND GND NM L=1.8e-07 W=2.2e-07 $X=182300 $Y=-148195 $D=0
M897 GND 76 383 GND NM L=1.8e-07 W=2.2e-07 $X=185960 $Y=-148195 $D=0
M898 1261 384 1252 GND NM L=1.8e-07 W=4.4e-07 $X=186000 $Y=-139615 $D=0
M899 386 383 GND GND NM L=1.8e-07 W=2.2e-07 $X=186760 $Y=-148195 $D=0
M900 1408 78 37 VDD PM L=1.8e-07 W=8.8e-07 $X=-167905 $Y=-98265 $D=4
M901 VDD 79 1408 VDD PM L=1.8e-07 W=8.8e-07 $X=-167475 $Y=-98265 $D=4
M902 1409 82 38 VDD PM L=1.8e-07 W=8.8e-07 $X=-156525 $Y=-98265 $D=4
M903 VDD 83 1409 VDD PM L=1.8e-07 W=8.8e-07 $X=-156095 $Y=-98265 $D=4
M904 1410 86 41 VDD PM L=1.8e-07 W=8.8e-07 $X=-145145 $Y=-98265 $D=4
M905 VDD 87 1410 VDD PM L=1.8e-07 W=8.8e-07 $X=-144715 $Y=-98265 $D=4
M906 1411 90 42 VDD PM L=1.8e-07 W=8.8e-07 $X=-133765 $Y=-98265 $D=4
M907 VDD 91 1411 VDD PM L=1.8e-07 W=8.8e-07 $X=-133335 $Y=-98265 $D=4
M908 1412 94 45 VDD PM L=1.8e-07 W=8.8e-07 $X=-122385 $Y=-98265 $D=4
M909 VDD 95 1412 VDD PM L=1.8e-07 W=8.8e-07 $X=-121955 $Y=-98265 $D=4
M910 1413 98 47 VDD PM L=1.8e-07 W=8.8e-07 $X=-111005 $Y=-98265 $D=4
M911 VDD 99 1413 VDD PM L=1.8e-07 W=8.8e-07 $X=-110575 $Y=-98265 $D=4
M912 1414 102 49 VDD PM L=1.8e-07 W=8.8e-07 $X=-99625 $Y=-98265 $D=4
M913 VDD 103 1414 VDD PM L=1.8e-07 W=8.8e-07 $X=-99195 $Y=-98265 $D=4
M914 1415 106 52 VDD PM L=1.8e-07 W=8.8e-07 $X=-88245 $Y=-98265 $D=4
M915 VDD 107 1415 VDD PM L=1.8e-07 W=8.8e-07 $X=-87815 $Y=-98265 $D=4
M916 1416 110 56 VDD PM L=1.8e-07 W=8.8e-07 $X=-76865 $Y=-98265 $D=4
M917 VDD 111 1416 VDD PM L=1.8e-07 W=8.8e-07 $X=-76435 $Y=-98265 $D=4
M918 1417 114 58 VDD PM L=1.8e-07 W=8.8e-07 $X=-65485 $Y=-98265 $D=4
M919 VDD 115 1417 VDD PM L=1.8e-07 W=8.8e-07 $X=-65055 $Y=-98265 $D=4
M920 1418 118 62 VDD PM L=1.8e-07 W=8.8e-07 $X=-54105 $Y=-98265 $D=4
M921 VDD 119 1418 VDD PM L=1.8e-07 W=8.8e-07 $X=-53675 $Y=-98265 $D=4
M922 1419 122 66 VDD PM L=1.8e-07 W=8.8e-07 $X=-42725 $Y=-98265 $D=4
M923 VDD 123 1419 VDD PM L=1.8e-07 W=8.8e-07 $X=-42295 $Y=-98265 $D=4
M924 1420 126 68 VDD PM L=1.8e-07 W=8.8e-07 $X=-31345 $Y=-98265 $D=4
M925 VDD 127 1420 VDD PM L=1.8e-07 W=8.8e-07 $X=-30915 $Y=-98265 $D=4
M926 1421 130 71 VDD PM L=1.8e-07 W=8.8e-07 $X=-19965 $Y=-98265 $D=4
M927 VDD 131 1421 VDD PM L=1.8e-07 W=8.8e-07 $X=-19535 $Y=-98265 $D=4
M928 1422 134 74 VDD PM L=1.8e-07 W=8.8e-07 $X=-8585 $Y=-98265 $D=4
M929 VDD 135 1422 VDD PM L=1.8e-07 W=8.8e-07 $X=-8155 $Y=-98265 $D=4
M930 1423 138 76 VDD PM L=1.8e-07 W=8.8e-07 $X=2795 $Y=-98265 $D=4
M931 VDD 140 1423 VDD PM L=1.8e-07 W=8.8e-07 $X=3225 $Y=-98265 $D=4
M932 406 6 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-55670 $D=4
M933 407 6 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-51170 $D=4
M934 408 6 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-49050 $D=4
M935 409 6 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-44550 $D=4
M936 VDD 414 144 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-42310 $D=4
M937 VDD 148 142 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-31720 $D=4
M938 157 153 142 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-29360 $D=4
M939 404 167 14 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=-5820 $D=4
M940 150 154 143 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=7130 $D=4
M941 VDD 149 143 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=9490 $D=4
M942 VDD 415 145 VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=20080 $D=4
M943 410 59 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=22320 $D=4
M944 411 59 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=26820 $D=4
M945 412 59 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=28940 $D=4
M946 413 59 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17440 $Y=33440 $D=4
M947 405 166 14 VDD PM L=1.8e-07 W=4.4e-07 $X=17480 $Y=-16410 $D=4
M948 414 146 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-42310 $D=4
M949 148 144 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-31720 $D=4
M950 148 151 157 VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=-29360 $D=4
M951 149 152 150 VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=7130 $D=4
M952 149 145 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=9490 $D=4
M953 415 147 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18160 $Y=20080 $D=4
M954 VDD 417 404 VDD PM L=1.8e-07 W=8.8e-07 $X=18200 $Y=-6260 $D=4
M955 VDD 416 405 VDD PM L=1.8e-07 W=8.8e-07 $X=18240 $Y=-16410 $D=4
M956 VDD 160 414 VDD PM L=1.8e-07 W=4.4e-07 $X=18880 $Y=-42310 $D=4
M957 VDD 155 148 VDD PM L=1.8e-07 W=4.4e-07 $X=18880 $Y=-31720 $D=4
M958 VDD 156 149 VDD PM L=1.8e-07 W=4.4e-07 $X=18880 $Y=9490 $D=4
M959 VDD 161 415 VDD PM L=1.8e-07 W=4.4e-07 $X=18880 $Y=20080 $D=4
M960 1424 157 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=18960 $Y=-16410 $D=4
M961 417 150 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=18960 $Y=-5820 $D=4
M962 416 150 1424 VDD PM L=1.8e-07 W=8.8e-07 $X=19390 $Y=-16410 $D=4
M963 155 406 11 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-55550 $D=4
M964 146 407 9 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-51070 $D=4
M965 188 408 7 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-48930 $D=4
M966 205 409 8 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=-44450 $D=4
M967 207 410 65 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=22440 $D=4
M968 189 411 63 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=26920 $D=4
M969 147 412 73 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=29060 $D=4
M970 156 413 70 VDD PM L=1.8e-07 W=2.2e-07 $X=19460 $Y=33540 $D=4
M971 VDD 157 417 VDD PM L=1.8e-07 W=4.4e-07 $X=19680 $Y=-5820 $D=4
M972 420 177 151 VDD PM L=1.8e-07 W=4.4e-07 $X=20100 $Y=-29360 $D=4
M973 421 178 152 VDD PM L=1.8e-07 W=4.4e-07 $X=20100 $Y=7130 $D=4
M974 418 173 151 VDD PM L=1.8e-07 W=4.4e-07 $X=20150 $Y=-18770 $D=4
M975 419 174 152 VDD PM L=1.8e-07 W=4.4e-07 $X=20150 $Y=-3460 $D=4
M976 GND 6 155 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-55550 $D=4
M977 GND 6 146 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-51070 $D=4
M978 GND 6 188 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-48930 $D=4
M979 GND 6 205 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=-44450 $D=4
M980 GND 59 207 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=22440 $D=4
M981 GND 59 189 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=26920 $D=4
M982 GND 59 147 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=29060 $D=4
M983 GND 59 156 VDD PM L=1.8e-07 W=2.2e-07 $X=20260 $Y=33540 $D=4
M984 422 414 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20820 $Y=-42310 $D=4
M985 423 148 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20820 $Y=-31720 $D=4
M986 424 149 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20820 $Y=9490 $D=4
M987 425 415 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=20820 $Y=20080 $D=4
M988 VDD 157 432 VDD PM L=1.8e-07 W=8.8e-07 $X=21330 $Y=-16410 $D=4
M989 1425 146 422 VDD PM L=1.8e-07 W=8.8e-07 $X=21580 $Y=-42310 $D=4
M990 1426 144 423 VDD PM L=1.8e-07 W=8.8e-07 $X=21580 $Y=-32160 $D=4
M991 1427 145 424 VDD PM L=1.8e-07 W=8.8e-07 $X=21580 $Y=9490 $D=4
M992 1428 147 425 VDD PM L=1.8e-07 W=8.8e-07 $X=21580 $Y=19640 $D=4
M993 426 417 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=21620 $Y=-5820 $D=4
M994 VDD 160 1425 VDD PM L=1.8e-07 W=8.8e-07 $X=22010 $Y=-42310 $D=4
M995 VDD 155 1426 VDD PM L=1.8e-07 W=8.8e-07 $X=22010 $Y=-32160 $D=4
M996 VDD 156 1427 VDD PM L=1.8e-07 W=8.8e-07 $X=22010 $Y=9490 $D=4
M997 VDD 161 1428 VDD PM L=1.8e-07 W=8.8e-07 $X=22010 $Y=19640 $D=4
M998 431 177 153 VDD PM L=1.8e-07 W=4.4e-07 $X=22050 $Y=-29360 $D=4
M999 432 150 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=22050 $Y=-16410 $D=4
M1000 433 178 154 VDD PM L=1.8e-07 W=4.4e-07 $X=22050 $Y=7130 $D=4
M1001 434 173 153 VDD PM L=1.8e-07 W=4.4e-07 $X=22090 $Y=-18770 $D=4
M1002 435 174 154 VDD PM L=1.8e-07 W=4.4e-07 $X=22090 $Y=-3460 $D=4
M1003 436 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=-55670 $D=4
M1004 437 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=-51170 $D=4
M1005 438 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=-49050 $D=4
M1006 439 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=-44550 $D=4
M1007 440 61 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=22320 $D=4
M1008 441 61 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=26820 $D=4
M1009 442 61 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=28940 $D=4
M1010 443 61 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22290 $Y=33440 $D=4
M1011 1429 150 426 VDD PM L=1.8e-07 W=8.8e-07 $X=22380 $Y=-6260 $D=4
M1012 445 416 432 VDD PM L=1.8e-07 W=8.8e-07 $X=22770 $Y=-16410 $D=4
M1013 VDD 420 431 VDD PM L=1.8e-07 W=8.8e-07 $X=22810 $Y=-29360 $D=4
M1014 VDD 157 1429 VDD PM L=1.8e-07 W=8.8e-07 $X=22810 $Y=-6260 $D=4
M1015 VDD 421 433 VDD PM L=1.8e-07 W=8.8e-07 $X=22810 $Y=6690 $D=4
M1016 VDD 418 434 VDD PM L=1.8e-07 W=8.8e-07 $X=22850 $Y=-19210 $D=4
M1017 VDD 419 435 VDD PM L=1.8e-07 W=8.8e-07 $X=22850 $Y=-3460 $D=4
M1018 420 158 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23570 $Y=-29360 $D=4
M1019 1430 162 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=23570 $Y=-19210 $D=4
M1020 1431 163 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=23570 $Y=-3460 $D=4
M1021 421 159 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23570 $Y=7130 $D=4
M1022 170 422 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23950 $Y=-42310 $D=4
M1023 158 423 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23950 $Y=-31720 $D=4
M1024 159 424 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23950 $Y=9490 $D=4
M1025 171 425 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=23950 $Y=20080 $D=4
M1026 418 158 1430 VDD PM L=1.8e-07 W=8.8e-07 $X=24000 $Y=-19210 $D=4
M1027 419 159 1431 VDD PM L=1.8e-07 W=8.8e-07 $X=24000 $Y=-3460 $D=4
M1028 VDD 162 420 VDD PM L=1.8e-07 W=4.4e-07 $X=24290 $Y=-29360 $D=4
M1029 VDD 163 421 VDD PM L=1.8e-07 W=4.4e-07 $X=24290 $Y=7130 $D=4
M1030 160 436 11 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-55550 $D=4
M1031 186 437 9 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-51070 $D=4
M1032 213 438 7 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-48930 $D=4
M1033 235 439 8 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=-44450 $D=4
M1034 236 440 65 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=22440 $D=4
M1035 214 441 63 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=26920 $D=4
M1036 187 442 73 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=29060 $D=4
M1037 161 443 70 VDD PM L=1.8e-07 W=2.2e-07 $X=24310 $Y=33540 $D=4
M1038 446 445 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=24710 $Y=-16410 $D=4
M1039 447 426 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=24750 $Y=-6260 $D=4
M1040 GND 10 160 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-55550 $D=4
M1041 GND 10 186 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-51070 $D=4
M1042 GND 10 213 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-48930 $D=4
M1043 GND 10 235 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=-44450 $D=4
M1044 GND 61 236 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=22440 $D=4
M1045 GND 61 214 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=26920 $D=4
M1046 GND 61 187 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=29060 $D=4
M1047 GND 61 161 VDD PM L=1.8e-07 W=2.2e-07 $X=25110 $Y=33540 $D=4
M1048 16 166 446 VDD PM L=1.8e-07 W=4.4e-07 $X=25470 $Y=-16410 $D=4
M1049 16 167 447 VDD PM L=1.8e-07 W=4.4e-07 $X=25510 $Y=-5820 $D=4
M1050 VDD 486 164 VDD PM L=1.8e-07 W=8.8e-07 $X=25930 $Y=-42310 $D=4
M1051 VDD 487 165 VDD PM L=1.8e-07 W=8.8e-07 $X=25930 $Y=19640 $D=4
M1052 VDD 162 451 VDD PM L=1.8e-07 W=8.8e-07 $X=25940 $Y=-19210 $D=4
M1053 VDD 163 452 VDD PM L=1.8e-07 W=8.8e-07 $X=25940 $Y=-3460 $D=4
M1054 VDD 456 162 VDD PM L=1.8e-07 W=4.4e-07 $X=26010 $Y=-31720 $D=4
M1055 VDD 457 163 VDD PM L=1.8e-07 W=4.4e-07 $X=26010 $Y=9490 $D=4
M1056 449 420 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=26230 $Y=-29360 $D=4
M1057 450 421 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=26230 $Y=7130 $D=4
M1058 451 158 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=26660 $Y=-19210 $D=4
M1059 452 159 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=26660 $Y=-3460 $D=4
M1060 456 164 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=26730 $Y=-31720 $D=4
M1061 457 165 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=26730 $Y=9490 $D=4
M1062 1432 158 449 VDD PM L=1.8e-07 W=8.8e-07 $X=26990 $Y=-29360 $D=4
M1063 1433 159 450 VDD PM L=1.8e-07 W=8.8e-07 $X=26990 $Y=6690 $D=4
M1064 458 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=-55670 $D=4
M1065 459 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=-51170 $D=4
M1066 460 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=-49050 $D=4
M1067 461 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=-44550 $D=4
M1068 462 53 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=22320 $D=4
M1069 463 53 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=26820 $D=4
M1070 464 53 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=28940 $D=4
M1071 465 53 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=27140 $Y=33440 $D=4
M1072 466 418 451 VDD PM L=1.8e-07 W=8.8e-07 $X=27380 $Y=-19210 $D=4
M1073 467 419 452 VDD PM L=1.8e-07 W=8.8e-07 $X=27380 $Y=-3460 $D=4
M1074 VDD 162 1432 VDD PM L=1.8e-07 W=8.8e-07 $X=27420 $Y=-29360 $D=4
M1075 VDD 163 1433 VDD PM L=1.8e-07 W=8.8e-07 $X=27420 $Y=6690 $D=4
M1076 VDD 170 456 VDD PM L=1.8e-07 W=4.4e-07 $X=27450 $Y=-31720 $D=4
M1077 VDD 171 457 VDD PM L=1.8e-07 W=4.4e-07 $X=27450 $Y=9490 $D=4
M1078 469 193 166 VDD PM L=1.8e-07 W=4.4e-07 $X=27560 $Y=-5820 $D=4
M1079 468 190 166 VDD PM L=1.8e-07 W=4.4e-07 $X=27610 $Y=-16410 $D=4
M1080 VDD 188 479 VDD PM L=1.8e-07 W=8.8e-07 $X=27870 $Y=-42310 $D=4
M1081 VDD 189 482 VDD PM L=1.8e-07 W=8.8e-07 $X=27870 $Y=19640 $D=4
M1082 1434 188 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=28590 $Y=-42310 $D=4
M1083 1435 189 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=28590 $Y=19640 $D=4
M1084 486 186 1434 VDD PM L=1.8e-07 W=8.8e-07 $X=29020 $Y=-42310 $D=4
M1085 487 187 1435 VDD PM L=1.8e-07 W=8.8e-07 $X=29020 $Y=19640 $D=4
M1086 175 458 11 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-55550 $D=4
M1087 182 459 9 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-51070 $D=4
M1088 168 460 7 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-48930 $D=4
M1089 244 461 8 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=-44450 $D=4
M1090 245 462 65 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=22440 $D=4
M1091 169 463 63 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=26920 $D=4
M1092 183 464 73 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=29060 $D=4
M1093 176 465 70 VDD PM L=1.8e-07 W=2.2e-07 $X=29160 $Y=33540 $D=4
M1094 471 466 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=29320 $Y=-19210 $D=4
M1095 472 467 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=29320 $Y=-3460 $D=4
M1096 473 449 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=29360 $Y=-29360 $D=4
M1097 474 450 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=29360 $Y=6690 $D=4
M1098 477 456 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29390 $Y=-31720 $D=4
M1099 478 457 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29390 $Y=9490 $D=4
M1100 475 193 167 VDD PM L=1.8e-07 W=4.4e-07 $X=29510 $Y=-5820 $D=4
M1101 476 190 167 VDD PM L=1.8e-07 W=4.4e-07 $X=29550 $Y=-16410 $D=4
M1102 479 175 486 VDD PM L=1.8e-07 W=8.8e-07 $X=29740 $Y=-42310 $D=4
M1103 482 176 487 VDD PM L=1.8e-07 W=8.8e-07 $X=29740 $Y=19640 $D=4
M1104 GND 12 175 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-55550 $D=4
M1105 GND 12 182 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-51070 $D=4
M1106 GND 12 168 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-48930 $D=4
M1107 GND 12 244 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=-44450 $D=4
M1108 GND 53 245 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=22440 $D=4
M1109 GND 53 169 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=26920 $D=4
M1110 GND 53 183 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=29060 $D=4
M1111 GND 53 176 VDD PM L=1.8e-07 W=2.2e-07 $X=29960 $Y=33540 $D=4
M1112 181 173 471 VDD PM L=1.8e-07 W=4.4e-07 $X=30080 $Y=-18770 $D=4
M1113 172 174 472 VDD PM L=1.8e-07 W=4.4e-07 $X=30080 $Y=-3460 $D=4
M1114 181 177 473 VDD PM L=1.8e-07 W=4.4e-07 $X=30120 $Y=-29360 $D=4
M1115 172 178 474 VDD PM L=1.8e-07 W=4.4e-07 $X=30120 $Y=7130 $D=4
M1116 1436 164 477 VDD PM L=1.8e-07 W=8.8e-07 $X=30150 $Y=-32160 $D=4
M1117 1437 165 478 VDD PM L=1.8e-07 W=8.8e-07 $X=30150 $Y=9490 $D=4
M1118 VDD 469 475 VDD PM L=1.8e-07 W=8.8e-07 $X=30270 $Y=-6260 $D=4
M1119 VDD 468 476 VDD PM L=1.8e-07 W=8.8e-07 $X=30310 $Y=-16410 $D=4
M1120 VDD 186 479 VDD PM L=1.8e-07 W=8.8e-07 $X=30460 $Y=-42310 $D=4
M1121 VDD 187 482 VDD PM L=1.8e-07 W=8.8e-07 $X=30460 $Y=19640 $D=4
M1122 VDD 170 1436 VDD PM L=1.8e-07 W=8.8e-07 $X=30580 $Y=-32160 $D=4
M1123 VDD 171 1437 VDD PM L=1.8e-07 W=8.8e-07 $X=30580 $Y=9490 $D=4
M1124 1438 181 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=31030 $Y=-16410 $D=4
M1125 469 172 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31030 $Y=-5820 $D=4
M1126 1439 186 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=31180 $Y=-42310 $D=4
M1127 1440 187 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=31180 $Y=19640 $D=4
M1128 468 172 1438 VDD PM L=1.8e-07 W=8.8e-07 $X=31460 $Y=-16410 $D=4
M1129 1441 188 1439 VDD PM L=1.8e-07 W=8.8e-07 $X=31610 $Y=-42310 $D=4
M1130 1442 189 1440 VDD PM L=1.8e-07 W=8.8e-07 $X=31610 $Y=19640 $D=4
M1131 VDD 181 469 VDD PM L=1.8e-07 W=4.4e-07 $X=31750 $Y=-5820 $D=4
M1132 488 13 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=-55670 $D=4
M1133 489 13 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=-51170 $D=4
M1134 490 13 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=-49050 $D=4
M1135 491 13 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=-44550 $D=4
M1136 492 54 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=22320 $D=4
M1137 493 54 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=26820 $D=4
M1138 494 54 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=28940 $D=4
M1139 495 54 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31990 $Y=33440 $D=4
M1140 513 175 1441 VDD PM L=1.8e-07 W=8.8e-07 $X=32040 $Y=-42310 $D=4
M1141 514 176 1442 VDD PM L=1.8e-07 W=8.8e-07 $X=32040 $Y=19640 $D=4
M1142 498 203 173 VDD PM L=1.8e-07 W=4.4e-07 $X=32170 $Y=-29360 $D=4
M1143 499 204 174 VDD PM L=1.8e-07 W=4.4e-07 $X=32170 $Y=7130 $D=4
M1144 496 199 173 VDD PM L=1.8e-07 W=4.4e-07 $X=32220 $Y=-18770 $D=4
M1145 497 200 174 VDD PM L=1.8e-07 W=4.4e-07 $X=32220 $Y=-3460 $D=4
M1146 184 477 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=32520 $Y=-31720 $D=4
M1147 185 478 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=32520 $Y=9490 $D=4
M1148 505 486 513 VDD PM L=1.8e-07 W=8.8e-07 $X=32760 $Y=-42310 $D=4
M1149 508 487 514 VDD PM L=1.8e-07 W=8.8e-07 $X=32760 $Y=19640 $D=4
M1150 VDD 181 503 VDD PM L=1.8e-07 W=8.8e-07 $X=33400 $Y=-16410 $D=4
M1151 VDD 175 505 VDD PM L=1.8e-07 W=8.8e-07 $X=33480 $Y=-42310 $D=4
M1152 VDD 176 508 VDD PM L=1.8e-07 W=8.8e-07 $X=33480 $Y=19640 $D=4
M1153 501 469 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=33690 $Y=-5820 $D=4
M1154 179 488 11 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-55550 $D=4
M1155 232 489 9 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-51070 $D=4
M1156 250 490 7 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-48930 $D=4
M1157 278 491 8 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=-44450 $D=4
M1158 283 492 65 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=22440 $D=4
M1159 251 493 63 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=26920 $D=4
M1160 233 494 73 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=29060 $D=4
M1161 180 495 70 VDD PM L=1.8e-07 W=2.2e-07 $X=34010 $Y=33540 $D=4
M1162 502 203 177 VDD PM L=1.8e-07 W=4.4e-07 $X=34120 $Y=-29360 $D=4
M1163 503 172 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=34120 $Y=-16410 $D=4
M1164 504 204 178 VDD PM L=1.8e-07 W=4.4e-07 $X=34120 $Y=7130 $D=4
M1165 509 199 177 VDD PM L=1.8e-07 W=4.4e-07 $X=34160 $Y=-18770 $D=4
M1166 510 200 178 VDD PM L=1.8e-07 W=4.4e-07 $X=34160 $Y=-3460 $D=4
M1167 505 188 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=34200 $Y=-42310 $D=4
M1168 508 189 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=34200 $Y=19640 $D=4
M1169 1443 172 501 VDD PM L=1.8e-07 W=8.8e-07 $X=34450 $Y=-6260 $D=4
M1170 VDD 537 191 VDD PM L=1.8e-07 W=8.8e-07 $X=34500 $Y=-32160 $D=4
M1171 VDD 538 192 VDD PM L=1.8e-07 W=8.8e-07 $X=34500 $Y=9490 $D=4
M1172 GND 13 179 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-55550 $D=4
M1173 GND 13 232 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-51070 $D=4
M1174 GND 13 250 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-48930 $D=4
M1175 GND 13 278 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=-44450 $D=4
M1176 GND 54 283 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=22440 $D=4
M1177 GND 54 251 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=26920 $D=4
M1178 GND 54 233 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=29060 $D=4
M1179 GND 54 180 VDD PM L=1.8e-07 W=2.2e-07 $X=34810 $Y=33540 $D=4
M1180 515 468 503 VDD PM L=1.8e-07 W=8.8e-07 $X=34840 $Y=-16410 $D=4
M1181 VDD 498 502 VDD PM L=1.8e-07 W=8.8e-07 $X=34880 $Y=-29360 $D=4
M1182 VDD 181 1443 VDD PM L=1.8e-07 W=8.8e-07 $X=34880 $Y=-6260 $D=4
M1183 VDD 499 504 VDD PM L=1.8e-07 W=8.8e-07 $X=34880 $Y=6690 $D=4
M1184 VDD 186 505 VDD PM L=1.8e-07 W=8.8e-07 $X=34920 $Y=-42310 $D=4
M1185 VDD 496 509 VDD PM L=1.8e-07 W=8.8e-07 $X=34920 $Y=-19210 $D=4
M1186 VDD 497 510 VDD PM L=1.8e-07 W=8.8e-07 $X=34920 $Y=-3460 $D=4
M1187 VDD 187 508 VDD PM L=1.8e-07 W=8.8e-07 $X=34920 $Y=19640 $D=4
M1188 194 513 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35640 $Y=-42310 $D=4
M1189 498 184 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=35640 $Y=-29360 $D=4
M1190 1444 191 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35640 $Y=-19210 $D=4
M1191 1445 192 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35640 $Y=-3460 $D=4
M1192 499 185 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=35640 $Y=7130 $D=4
M1193 195 514 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35640 $Y=19640 $D=4
M1194 496 184 1444 VDD PM L=1.8e-07 W=8.8e-07 $X=36070 $Y=-19210 $D=4
M1195 497 185 1445 VDD PM L=1.8e-07 W=8.8e-07 $X=36070 $Y=-3460 $D=4
M1196 VDD 191 498 VDD PM L=1.8e-07 W=4.4e-07 $X=36360 $Y=-29360 $D=4
M1197 VDD 192 499 VDD PM L=1.8e-07 W=4.4e-07 $X=36360 $Y=7130 $D=4
M1198 VDD 197 520 VDD PM L=1.8e-07 W=8.8e-07 $X=36440 $Y=-32160 $D=4
M1199 VDD 198 521 VDD PM L=1.8e-07 W=8.8e-07 $X=36440 $Y=9490 $D=4
M1200 517 515 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=36780 $Y=-16410 $D=4
M1201 518 501 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=36820 $Y=-6260 $D=4
M1202 1446 197 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=37160 $Y=-32160 $D=4
M1203 1447 198 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=37160 $Y=9490 $D=4
M1204 18 190 517 VDD PM L=1.8e-07 W=4.4e-07 $X=37540 $Y=-16410 $D=4
M1205 18 193 518 VDD PM L=1.8e-07 W=4.4e-07 $X=37580 $Y=-5820 $D=4
M1206 537 201 1446 VDD PM L=1.8e-07 W=8.8e-07 $X=37590 $Y=-32160 $D=4
M1207 538 202 1447 VDD PM L=1.8e-07 W=8.8e-07 $X=37590 $Y=9490 $D=4
M1208 VDD 528 201 VDD PM L=1.8e-07 W=4.4e-07 $X=37660 $Y=-42310 $D=4
M1209 VDD 529 202 VDD PM L=1.8e-07 W=4.4e-07 $X=37660 $Y=20080 $D=4
M1210 VDD 191 526 VDD PM L=1.8e-07 W=8.8e-07 $X=38010 $Y=-19210 $D=4
M1211 VDD 192 527 VDD PM L=1.8e-07 W=8.8e-07 $X=38010 $Y=-3460 $D=4
M1212 524 498 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=38300 $Y=-29360 $D=4
M1213 525 499 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=38300 $Y=7130 $D=4
M1214 520 194 537 VDD PM L=1.8e-07 W=8.8e-07 $X=38310 $Y=-32160 $D=4
M1215 521 195 538 VDD PM L=1.8e-07 W=8.8e-07 $X=38310 $Y=9490 $D=4
M1216 528 182 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=38380 $Y=-42310 $D=4
M1217 529 183 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=38380 $Y=20080 $D=4
M1218 526 184 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=38730 $Y=-19210 $D=4
M1219 527 185 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=38730 $Y=-3460 $D=4
M1220 VDD 201 520 VDD PM L=1.8e-07 W=8.8e-07 $X=39030 $Y=-32160 $D=4
M1221 VDD 202 521 VDD PM L=1.8e-07 W=8.8e-07 $X=39030 $Y=9490 $D=4
M1222 1448 184 524 VDD PM L=1.8e-07 W=8.8e-07 $X=39060 $Y=-29360 $D=4
M1223 1449 185 525 VDD PM L=1.8e-07 W=8.8e-07 $X=39060 $Y=6690 $D=4
M1224 VDD 179 528 VDD PM L=1.8e-07 W=4.4e-07 $X=39100 $Y=-42310 $D=4
M1225 VDD 180 529 VDD PM L=1.8e-07 W=4.4e-07 $X=39100 $Y=20080 $D=4
M1226 532 496 526 VDD PM L=1.8e-07 W=8.8e-07 $X=39450 $Y=-19210 $D=4
M1227 533 497 527 VDD PM L=1.8e-07 W=8.8e-07 $X=39450 $Y=-3460 $D=4
M1228 VDD 191 1448 VDD PM L=1.8e-07 W=8.8e-07 $X=39490 $Y=-29360 $D=4
M1229 VDD 192 1449 VDD PM L=1.8e-07 W=8.8e-07 $X=39490 $Y=6690 $D=4
M1230 535 215 190 VDD PM L=1.8e-07 W=4.4e-07 $X=39630 $Y=-5820 $D=4
M1231 534 212 190 VDD PM L=1.8e-07 W=4.4e-07 $X=39680 $Y=-16410 $D=4
M1232 1450 201 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=39750 $Y=-32160 $D=4
M1233 1451 202 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=39750 $Y=9490 $D=4
M1234 1452 197 1450 VDD PM L=1.8e-07 W=8.8e-07 $X=40180 $Y=-32160 $D=4
M1235 1453 198 1451 VDD PM L=1.8e-07 W=8.8e-07 $X=40180 $Y=9490 $D=4
M1236 554 194 1452 VDD PM L=1.8e-07 W=8.8e-07 $X=40610 $Y=-32160 $D=4
M1237 555 195 1453 VDD PM L=1.8e-07 W=8.8e-07 $X=40610 $Y=9490 $D=4
M1238 539 528 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=41040 $Y=-42310 $D=4
M1239 540 529 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=41040 $Y=20080 $D=4
M1240 551 537 554 VDD PM L=1.8e-07 W=8.8e-07 $X=41330 $Y=-32160 $D=4
M1241 552 538 555 VDD PM L=1.8e-07 W=8.8e-07 $X=41330 $Y=9490 $D=4
M1242 541 532 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41390 $Y=-19210 $D=4
M1243 542 533 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41390 $Y=-3460 $D=4
M1244 543 524 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41430 $Y=-29360 $D=4
M1245 544 525 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41430 $Y=6690 $D=4
M1246 545 215 193 VDD PM L=1.8e-07 W=4.4e-07 $X=41580 $Y=-5820 $D=4
M1247 546 212 193 VDD PM L=1.8e-07 W=4.4e-07 $X=41620 $Y=-16410 $D=4
M1248 1454 182 539 VDD PM L=1.8e-07 W=8.8e-07 $X=41800 $Y=-42310 $D=4
M1249 1455 183 540 VDD PM L=1.8e-07 W=8.8e-07 $X=41800 $Y=19640 $D=4
M1250 VDD 194 551 VDD PM L=1.8e-07 W=8.8e-07 $X=42050 $Y=-32160 $D=4
M1251 VDD 195 552 VDD PM L=1.8e-07 W=8.8e-07 $X=42050 $Y=9490 $D=4
M1252 206 199 541 VDD PM L=1.8e-07 W=4.4e-07 $X=42150 $Y=-18770 $D=4
M1253 196 200 542 VDD PM L=1.8e-07 W=4.4e-07 $X=42150 $Y=-3460 $D=4
M1254 206 203 543 VDD PM L=1.8e-07 W=4.4e-07 $X=42190 $Y=-29360 $D=4
M1255 196 204 544 VDD PM L=1.8e-07 W=4.4e-07 $X=42190 $Y=7130 $D=4
M1256 VDD 179 1454 VDD PM L=1.8e-07 W=8.8e-07 $X=42230 $Y=-42310 $D=4
M1257 VDD 180 1455 VDD PM L=1.8e-07 W=8.8e-07 $X=42230 $Y=19640 $D=4
M1258 VDD 535 545 VDD PM L=1.8e-07 W=8.8e-07 $X=42340 $Y=-6260 $D=4
M1259 VDD 534 546 VDD PM L=1.8e-07 W=8.8e-07 $X=42380 $Y=-16410 $D=4
M1260 551 197 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42770 $Y=-32160 $D=4
M1261 552 198 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42770 $Y=9490 $D=4
M1262 1456 206 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=43100 $Y=-16410 $D=4
M1263 535 196 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=43100 $Y=-5820 $D=4
M1264 VDD 201 551 VDD PM L=1.8e-07 W=8.8e-07 $X=43490 $Y=-32160 $D=4
M1265 VDD 202 552 VDD PM L=1.8e-07 W=8.8e-07 $X=43490 $Y=9490 $D=4
M1266 534 196 1456 VDD PM L=1.8e-07 W=8.8e-07 $X=43530 $Y=-16410 $D=4
M1267 VDD 206 535 VDD PM L=1.8e-07 W=4.4e-07 $X=43820 $Y=-5820 $D=4
M1268 220 539 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=44170 $Y=-42310 $D=4
M1269 221 540 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=44170 $Y=20080 $D=4
M1270 208 554 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44210 $Y=-32160 $D=4
M1271 209 555 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44210 $Y=9490 $D=4
M1272 559 563 199 VDD PM L=1.8e-07 W=4.4e-07 $X=44240 $Y=-29360 $D=4
M1273 560 564 200 VDD PM L=1.8e-07 W=4.4e-07 $X=44240 $Y=7130 $D=4
M1274 557 561 199 VDD PM L=1.8e-07 W=4.4e-07 $X=44290 $Y=-18770 $D=4
M1275 558 562 200 VDD PM L=1.8e-07 W=4.4e-07 $X=44290 $Y=-3460 $D=4
M1276 VDD 206 567 VDD PM L=1.8e-07 W=8.8e-07 $X=45470 $Y=-16410 $D=4
M1277 565 535 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=45760 $Y=-5820 $D=4
M1278 VDD 599 210 VDD PM L=1.8e-07 W=8.8e-07 $X=46150 $Y=-32160 $D=4
M1279 VDD 600 211 VDD PM L=1.8e-07 W=8.8e-07 $X=46150 $Y=9490 $D=4
M1280 566 563 203 VDD PM L=1.8e-07 W=4.4e-07 $X=46190 $Y=-29360 $D=4
M1281 567 196 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=46190 $Y=-16410 $D=4
M1282 568 564 204 VDD PM L=1.8e-07 W=4.4e-07 $X=46190 $Y=7130 $D=4
M1283 VDD 574 197 VDD PM L=1.8e-07 W=4.4e-07 $X=46230 $Y=-42310 $D=4
M1284 570 561 203 VDD PM L=1.8e-07 W=4.4e-07 $X=46230 $Y=-18770 $D=4
M1285 571 562 204 VDD PM L=1.8e-07 W=4.4e-07 $X=46230 $Y=-3460 $D=4
M1286 VDD 575 198 VDD PM L=1.8e-07 W=4.4e-07 $X=46230 $Y=20080 $D=4
M1287 1457 196 565 VDD PM L=1.8e-07 W=8.8e-07 $X=46520 $Y=-6260 $D=4
M1288 573 534 567 VDD PM L=1.8e-07 W=8.8e-07 $X=46910 $Y=-16410 $D=4
M1289 574 205 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=46950 $Y=-42310 $D=4
M1290 VDD 559 566 VDD PM L=1.8e-07 W=8.8e-07 $X=46950 $Y=-29360 $D=4
M1291 VDD 206 1457 VDD PM L=1.8e-07 W=8.8e-07 $X=46950 $Y=-6260 $D=4
M1292 VDD 560 568 VDD PM L=1.8e-07 W=8.8e-07 $X=46950 $Y=6690 $D=4
M1293 575 207 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=46950 $Y=20080 $D=4
M1294 VDD 557 570 VDD PM L=1.8e-07 W=8.8e-07 $X=46990 $Y=-19210 $D=4
M1295 VDD 558 571 VDD PM L=1.8e-07 W=8.8e-07 $X=46990 $Y=-3460 $D=4
M1296 VDD 213 574 VDD PM L=1.8e-07 W=4.4e-07 $X=47670 $Y=-42310 $D=4
M1297 VDD 214 575 VDD PM L=1.8e-07 W=4.4e-07 $X=47670 $Y=20080 $D=4
M1298 559 208 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=47710 $Y=-29360 $D=4
M1299 1458 210 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=47710 $Y=-19210 $D=4
M1300 1459 211 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=47710 $Y=-3460 $D=4
M1301 560 209 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=47710 $Y=7130 $D=4
M1302 VDD 218 582 VDD PM L=1.8e-07 W=8.8e-07 $X=48090 $Y=-32160 $D=4
M1303 VDD 219 583 VDD PM L=1.8e-07 W=8.8e-07 $X=48090 $Y=9490 $D=4
M1304 557 208 1458 VDD PM L=1.8e-07 W=8.8e-07 $X=48140 $Y=-19210 $D=4
M1305 558 209 1459 VDD PM L=1.8e-07 W=8.8e-07 $X=48140 $Y=-3460 $D=4
M1306 VDD 210 559 VDD PM L=1.8e-07 W=4.4e-07 $X=48430 $Y=-29360 $D=4
M1307 VDD 211 560 VDD PM L=1.8e-07 W=4.4e-07 $X=48430 $Y=7130 $D=4
M1308 1460 218 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48810 $Y=-32160 $D=4
M1309 1461 219 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48810 $Y=9490 $D=4
M1310 577 573 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48850 $Y=-16410 $D=4
M1311 578 565 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48890 $Y=-6260 $D=4
M1312 599 220 1460 VDD PM L=1.8e-07 W=8.8e-07 $X=49240 $Y=-32160 $D=4
M1313 600 221 1461 VDD PM L=1.8e-07 W=8.8e-07 $X=49240 $Y=9490 $D=4
M1314 579 574 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=49610 $Y=-42310 $D=4
M1315 29 212 577 VDD PM L=1.8e-07 W=4.4e-07 $X=49610 $Y=-16410 $D=4
M1316 580 575 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=49610 $Y=20080 $D=4
M1317 29 215 578 VDD PM L=1.8e-07 W=4.4e-07 $X=49650 $Y=-5820 $D=4
M1318 582 216 599 VDD PM L=1.8e-07 W=8.8e-07 $X=49960 $Y=-32160 $D=4
M1319 583 217 600 VDD PM L=1.8e-07 W=8.8e-07 $X=49960 $Y=9490 $D=4
M1320 VDD 210 590 VDD PM L=1.8e-07 W=8.8e-07 $X=50080 $Y=-19210 $D=4
M1321 VDD 211 591 VDD PM L=1.8e-07 W=8.8e-07 $X=50080 $Y=-3460 $D=4
M1322 1462 205 579 VDD PM L=1.8e-07 W=8.8e-07 $X=50370 $Y=-42310 $D=4
M1323 586 559 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=50370 $Y=-29360 $D=4
M1324 587 560 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=50370 $Y=7130 $D=4
M1325 1463 207 580 VDD PM L=1.8e-07 W=8.8e-07 $X=50370 $Y=19640 $D=4
M1326 VDD 220 582 VDD PM L=1.8e-07 W=8.8e-07 $X=50680 $Y=-32160 $D=4
M1327 VDD 221 583 VDD PM L=1.8e-07 W=8.8e-07 $X=50680 $Y=9490 $D=4
M1328 VDD 213 1462 VDD PM L=1.8e-07 W=8.8e-07 $X=50800 $Y=-42310 $D=4
M1329 590 208 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50800 $Y=-19210 $D=4
M1330 591 209 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50800 $Y=-3460 $D=4
M1331 VDD 214 1463 VDD PM L=1.8e-07 W=8.8e-07 $X=50800 $Y=19640 $D=4
M1332 1464 208 586 VDD PM L=1.8e-07 W=8.8e-07 $X=51130 $Y=-29360 $D=4
M1333 1465 209 587 VDD PM L=1.8e-07 W=8.8e-07 $X=51130 $Y=6690 $D=4
M1334 1466 220 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=51400 $Y=-32160 $D=4
M1335 1467 221 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=51400 $Y=9490 $D=4
M1336 594 557 590 VDD PM L=1.8e-07 W=8.8e-07 $X=51520 $Y=-19210 $D=4
M1337 595 558 591 VDD PM L=1.8e-07 W=8.8e-07 $X=51520 $Y=-3460 $D=4
M1338 VDD 210 1464 VDD PM L=1.8e-07 W=8.8e-07 $X=51560 $Y=-29360 $D=4
M1339 VDD 211 1465 VDD PM L=1.8e-07 W=8.8e-07 $X=51560 $Y=6690 $D=4
M1340 597 240 212 VDD PM L=1.8e-07 W=4.4e-07 $X=51700 $Y=-5820 $D=4
M1341 596 237 212 VDD PM L=1.8e-07 W=4.4e-07 $X=51750 $Y=-16410 $D=4
M1342 1468 218 1466 VDD PM L=1.8e-07 W=8.8e-07 $X=51830 $Y=-32160 $D=4
M1343 1469 219 1467 VDD PM L=1.8e-07 W=8.8e-07 $X=51830 $Y=9490 $D=4
M1344 612 216 1468 VDD PM L=1.8e-07 W=8.8e-07 $X=52260 $Y=-32160 $D=4
M1345 613 217 1469 VDD PM L=1.8e-07 W=8.8e-07 $X=52260 $Y=9490 $D=4
M1346 218 579 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=52740 $Y=-42310 $D=4
M1347 219 580 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=52740 $Y=20080 $D=4
M1348 609 599 612 VDD PM L=1.8e-07 W=8.8e-07 $X=52980 $Y=-32160 $D=4
M1349 610 600 613 VDD PM L=1.8e-07 W=8.8e-07 $X=52980 $Y=9490 $D=4
M1350 601 594 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53460 $Y=-19210 $D=4
M1351 602 595 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53460 $Y=-3460 $D=4
M1352 603 586 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53500 $Y=-29360 $D=4
M1353 604 587 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=53500 $Y=6690 $D=4
M1354 605 240 215 VDD PM L=1.8e-07 W=4.4e-07 $X=53650 $Y=-5820 $D=4
M1355 606 237 215 VDD PM L=1.8e-07 W=4.4e-07 $X=53690 $Y=-16410 $D=4
M1356 VDD 216 609 VDD PM L=1.8e-07 W=8.8e-07 $X=53700 $Y=-32160 $D=4
M1357 VDD 217 610 VDD PM L=1.8e-07 W=8.8e-07 $X=53700 $Y=9490 $D=4
M1358 225 561 601 VDD PM L=1.8e-07 W=4.4e-07 $X=54220 $Y=-18770 $D=4
M1359 222 562 602 VDD PM L=1.8e-07 W=4.4e-07 $X=54220 $Y=-3460 $D=4
M1360 225 563 603 VDD PM L=1.8e-07 W=4.4e-07 $X=54260 $Y=-29360 $D=4
M1361 222 564 604 VDD PM L=1.8e-07 W=4.4e-07 $X=54260 $Y=7130 $D=4
M1362 VDD 597 605 VDD PM L=1.8e-07 W=8.8e-07 $X=54410 $Y=-6260 $D=4
M1363 609 218 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54420 $Y=-32160 $D=4
M1364 610 219 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54420 $Y=9490 $D=4
M1365 VDD 596 606 VDD PM L=1.8e-07 W=8.8e-07 $X=54450 $Y=-16410 $D=4
M1366 VDD 639 216 VDD PM L=1.8e-07 W=8.8e-07 $X=54720 $Y=-42310 $D=4
M1367 VDD 640 217 VDD PM L=1.8e-07 W=8.8e-07 $X=54720 $Y=19640 $D=4
M1368 VDD 220 609 VDD PM L=1.8e-07 W=8.8e-07 $X=55140 $Y=-32160 $D=4
M1369 VDD 221 610 VDD PM L=1.8e-07 W=8.8e-07 $X=55140 $Y=9490 $D=4
M1370 1470 225 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=55170 $Y=-16410 $D=4
M1371 597 222 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=55170 $Y=-5820 $D=4
M1372 596 222 1470 VDD PM L=1.8e-07 W=8.8e-07 $X=55600 $Y=-16410 $D=4
M1373 229 612 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=55860 $Y=-32160 $D=4
M1374 230 613 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=55860 $Y=9490 $D=4
M1375 VDD 225 597 VDD PM L=1.8e-07 W=4.4e-07 $X=55890 $Y=-5820 $D=4
M1376 624 20 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=56240 $Y=-18770 $D=4
M1377 625 14 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=56240 $Y=-3460 $D=4
M1378 VDD 561 563 VDD PM L=1.8e-07 W=4.4e-07 $X=56280 $Y=-29360 $D=4
M1379 VDD 562 564 VDD PM L=1.8e-07 W=4.4e-07 $X=56280 $Y=7130 $D=4
M1380 VDD 235 620 VDD PM L=1.8e-07 W=8.8e-07 $X=56660 $Y=-42310 $D=4
M1381 VDD 236 623 VDD PM L=1.8e-07 W=8.8e-07 $X=56660 $Y=19640 $D=4
M1382 561 223 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=57000 $Y=-29360 $D=4
M1383 562 224 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=57000 $Y=7130 $D=4
M1384 1471 235 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=57380 $Y=-42310 $D=4
M1385 1472 236 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=57380 $Y=19640 $D=4
M1386 VDD 225 619 VDD PM L=1.8e-07 W=8.8e-07 $X=57540 $Y=-16410 $D=4
M1387 VDD 229 561 VDD PM L=1.8e-07 W=4.4e-07 $X=57720 $Y=-29360 $D=4
M1388 VDD 230 562 VDD PM L=1.8e-07 W=4.4e-07 $X=57720 $Y=7130 $D=4
M1389 639 168 1471 VDD PM L=1.8e-07 W=8.8e-07 $X=57810 $Y=-42310 $D=4
M1390 640 169 1472 VDD PM L=1.8e-07 W=8.8e-07 $X=57810 $Y=19640 $D=4
M1391 618 597 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=57830 $Y=-5820 $D=4
M1392 VDD 628 223 VDD PM L=1.8e-07 W=4.4e-07 $X=57880 $Y=-31720 $D=4
M1393 VDD 629 224 VDD PM L=1.8e-07 W=4.4e-07 $X=57880 $Y=9490 $D=4
M1394 1473 CLK 615 VDD PM L=1.8e-07 W=8.8e-07 $X=58180 $Y=-19210 $D=4
M1395 1474 CLK 616 VDD PM L=1.8e-07 W=8.8e-07 $X=58180 $Y=-3460 $D=4
M1396 619 222 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=58260 $Y=-16410 $D=4
M1397 620 232 639 VDD PM L=1.8e-07 W=8.8e-07 $X=58530 $Y=-42310 $D=4
M1398 623 233 640 VDD PM L=1.8e-07 W=8.8e-07 $X=58530 $Y=19640 $D=4
M1399 1475 222 618 VDD PM L=1.8e-07 W=8.8e-07 $X=58590 $Y=-6260 $D=4
M1400 628 242 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=58600 $Y=-31720 $D=4
M1401 629 243 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=58600 $Y=9490 $D=4
M1402 1476 RST 1473 VDD PM L=1.8e-07 W=8.8e-07 $X=58610 $Y=-19210 $D=4
M1403 1477 RST 1474 VDD PM L=1.8e-07 W=8.8e-07 $X=58610 $Y=-3460 $D=4
M1404 627 596 619 VDD PM L=1.8e-07 W=8.8e-07 $X=58980 $Y=-16410 $D=4
M1405 VDD 225 1475 VDD PM L=1.8e-07 W=8.8e-07 $X=59020 $Y=-6260 $D=4
M1406 VDD 624 1476 VDD PM L=1.8e-07 W=8.8e-07 $X=59040 $Y=-19210 $D=4
M1407 VDD 625 1477 VDD PM L=1.8e-07 W=8.8e-07 $X=59040 $Y=-3460 $D=4
M1408 VDD 168 620 VDD PM L=1.8e-07 W=8.8e-07 $X=59250 $Y=-42310 $D=4
M1409 VDD 169 623 VDD PM L=1.8e-07 W=8.8e-07 $X=59250 $Y=19640 $D=4
M1410 VDD 238 628 VDD PM L=1.8e-07 W=4.4e-07 $X=59320 $Y=-31720 $D=4
M1411 VDD 239 629 VDD PM L=1.8e-07 W=4.4e-07 $X=59320 $Y=9490 $D=4
M1412 631 561 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=59660 $Y=-29360 $D=4
M1413 632 562 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=59660 $Y=7130 $D=4
M1414 633 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=59760 $Y=-19210 $D=4
M1415 634 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=59760 $Y=-3460 $D=4
M1416 1478 168 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=59970 $Y=-42310 $D=4
M1417 1479 169 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=59970 $Y=19640 $D=4
M1418 1480 235 1478 VDD PM L=1.8e-07 W=8.8e-07 $X=60400 $Y=-42310 $D=4
M1419 1481 236 1479 VDD PM L=1.8e-07 W=8.8e-07 $X=60400 $Y=19640 $D=4
M1420 1482 223 631 VDD PM L=1.8e-07 W=8.8e-07 $X=60420 $Y=-29360 $D=4
M1421 1483 224 632 VDD PM L=1.8e-07 W=8.8e-07 $X=60420 $Y=6690 $D=4
M1422 652 232 1480 VDD PM L=1.8e-07 W=8.8e-07 $X=60830 $Y=-42310 $D=4
M1423 653 233 1481 VDD PM L=1.8e-07 W=8.8e-07 $X=60830 $Y=19640 $D=4
M1424 VDD 229 1482 VDD PM L=1.8e-07 W=8.8e-07 $X=60850 $Y=-29360 $D=4
M1425 VDD 230 1483 VDD PM L=1.8e-07 W=8.8e-07 $X=60850 $Y=6690 $D=4
M1426 637 627 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=60920 $Y=-16410 $D=4
M1427 638 618 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=60960 $Y=-6260 $D=4
M1428 641 628 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=61260 $Y=-31720 $D=4
M1429 642 629 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=61260 $Y=9490 $D=4
M1430 647 639 652 VDD PM L=1.8e-07 W=8.8e-07 $X=61550 $Y=-42310 $D=4
M1431 650 640 653 VDD PM L=1.8e-07 W=8.8e-07 $X=61550 $Y=19640 $D=4
M1432 32 237 637 VDD PM L=1.8e-07 W=4.4e-07 $X=61680 $Y=-16410 $D=4
M1433 32 240 638 VDD PM L=1.8e-07 W=4.4e-07 $X=61720 $Y=-5820 $D=4
M1434 1484 242 641 VDD PM L=1.8e-07 W=8.8e-07 $X=62020 $Y=-32160 $D=4
M1435 1485 243 642 VDD PM L=1.8e-07 W=8.8e-07 $X=62020 $Y=9490 $D=4
M1436 VDD 232 647 VDD PM L=1.8e-07 W=8.8e-07 $X=62270 $Y=-42310 $D=4
M1437 VDD 233 650 VDD PM L=1.8e-07 W=8.8e-07 $X=62270 $Y=19640 $D=4
M1438 VDD 238 1484 VDD PM L=1.8e-07 W=8.8e-07 $X=62450 $Y=-32160 $D=4
M1439 VDD 239 1485 VDD PM L=1.8e-07 W=8.8e-07 $X=62450 $Y=9490 $D=4
M1440 VDD 633 Q3 VDD PM L=1.8e-07 W=8.8e-07 $X=62460 $Y=-19210 $D=4
M1441 VDD 634 Q8 VDD PM L=1.8e-07 W=8.8e-07 $X=62460 $Y=-3460 $D=4
M1442 252 631 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=62790 $Y=-29360 $D=4
M1443 246 632 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=62790 $Y=7130 $D=4
M1444 647 235 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=62990 $Y=-42310 $D=4
M1445 650 236 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=62990 $Y=19640 $D=4
M1446 VDD 168 647 VDD PM L=1.8e-07 W=8.8e-07 $X=63710 $Y=-42310 $D=4
M1447 VDD 169 650 VDD PM L=1.8e-07 W=8.8e-07 $X=63710 $Y=19640 $D=4
M1448 655 260 237 VDD PM L=1.8e-07 W=4.4e-07 $X=63770 $Y=-5820 $D=4
M1449 654 258 237 VDD PM L=1.8e-07 W=4.4e-07 $X=63820 $Y=-16410 $D=4
M1450 272 641 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=64390 $Y=-31720 $D=4
M1451 263 642 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=64390 $Y=9490 $D=4
M1452 238 652 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=64430 $Y=-42310 $D=4
M1453 239 653 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=64430 $Y=19640 $D=4
M1454 664 30 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=65160 $Y=-18770 $D=4
M1455 665 16 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=65160 $Y=-3460 $D=4
M1456 658 260 240 VDD PM L=1.8e-07 W=4.4e-07 $X=65720 $Y=-5820 $D=4
M1457 659 258 240 VDD PM L=1.8e-07 W=4.4e-07 $X=65760 $Y=-16410 $D=4
M1458 VDD 666 242 VDD PM L=1.8e-07 W=4.4e-07 $X=66450 $Y=-42310 $D=4
M1459 VDD 667 243 VDD PM L=1.8e-07 W=4.4e-07 $X=66450 $Y=20080 $D=4
M1460 VDD 655 658 VDD PM L=1.8e-07 W=8.8e-07 $X=66480 $Y=-6260 $D=4
M1461 VDD 654 659 VDD PM L=1.8e-07 W=8.8e-07 $X=66520 $Y=-16410 $D=4
M1462 1486 231 247 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-122795 $D=4
M1463 VDD 234 1487 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-121935 $D=4
M1464 1488 231 253 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-119175 $D=4
M1465 1489 241 1488 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-118745 $D=4
M1466 VDD ADD0 1489 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-118315 $D=4
M1467 1490 231 254 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-115555 $D=4
M1468 1491 ADD1 1490 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-115125 $D=4
M1469 VDD 234 1491 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-114695 $D=4
M1470 VDD ADD0 1492 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-111075 $D=4
M1471 1494 ADD1 1493 VDD PM L=1.8e-07 W=1.32e-06 $X=66940 $Y=-100645 $D=4
M1472 1495 CLK 661 VDD PM L=1.8e-07 W=8.8e-07 $X=67100 $Y=-19210 $D=4
M1473 1496 CLK 662 VDD PM L=1.8e-07 W=8.8e-07 $X=67100 $Y=-3460 $D=4
M1474 666 244 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=67170 $Y=-42310 $D=4
M1475 667 245 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=67170 $Y=20080 $D=4
M1476 1497 252 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=67240 $Y=-16410 $D=4
M1477 655 246 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=67240 $Y=-5820 $D=4
M1478 1498 RST 1495 VDD PM L=1.8e-07 W=8.8e-07 $X=67530 $Y=-19210 $D=4
M1479 1499 RST 1496 VDD PM L=1.8e-07 W=8.8e-07 $X=67530 $Y=-3460 $D=4
M1480 654 246 1497 VDD PM L=1.8e-07 W=8.8e-07 $X=67670 $Y=-16410 $D=4
M1481 VDD 250 666 VDD PM L=1.8e-07 W=4.4e-07 $X=67890 $Y=-42310 $D=4
M1482 VDD 251 667 VDD PM L=1.8e-07 W=4.4e-07 $X=67890 $Y=20080 $D=4
M1483 VDD 664 1498 VDD PM L=1.8e-07 W=8.8e-07 $X=67960 $Y=-19210 $D=4
M1484 VDD 252 655 VDD PM L=1.8e-07 W=4.4e-07 $X=67960 $Y=-5820 $D=4
M1485 VDD 665 1499 VDD PM L=1.8e-07 W=8.8e-07 $X=67960 $Y=-3460 $D=4
M1486 670 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=68680 $Y=-19210 $D=4
M1487 671 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=68680 $Y=-3460 $D=4
M1488 VDD 252 676 VDD PM L=1.8e-07 W=8.8e-07 $X=69610 $Y=-16410 $D=4
M1489 687 247 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-129795 $D=4
M1490 688 253 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-125155 $D=4
M1491 689 254 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-120515 $D=4
M1492 690 255 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-115875 $D=4
M1493 691 256 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-111235 $D=4
M1494 VDD 692 23 VDD PM L=1.8e-07 W=4.4e-07 $X=69740 $Y=-108535 $D=4
M1495 692 257 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-106595 $D=4
M1496 VDD 693 22 VDD PM L=1.8e-07 W=4.4e-07 $X=69740 $Y=-103895 $D=4
M1497 693 248 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-101955 $D=4
M1498 VDD CLK 693 VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-101235 $D=4
M1499 694 249 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-97315 $D=4
M1500 VDD CLK 694 VDD PM L=1.8e-07 W=8.8e-07 $X=69740 $Y=-96595 $D=4
M1501 673 666 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=69830 $Y=-42310 $D=4
M1502 674 667 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=69830 $Y=20080 $D=4
M1503 675 655 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=69900 $Y=-5820 $D=4
M1504 676 246 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=70330 $Y=-16410 $D=4
M1505 1500 244 673 VDD PM L=1.8e-07 W=8.8e-07 $X=70590 $Y=-42310 $D=4
M1506 1501 245 674 VDD PM L=1.8e-07 W=8.8e-07 $X=70590 $Y=19640 $D=4
M1507 1502 246 675 VDD PM L=1.8e-07 W=8.8e-07 $X=70660 $Y=-6260 $D=4
M1508 VDD 250 1500 VDD PM L=1.8e-07 W=8.8e-07 $X=71020 $Y=-42310 $D=4
M1509 VDD 251 1501 VDD PM L=1.8e-07 W=8.8e-07 $X=71020 $Y=19640 $D=4
M1510 680 654 676 VDD PM L=1.8e-07 W=8.8e-07 $X=71050 $Y=-16410 $D=4
M1511 VDD 252 1502 VDD PM L=1.8e-07 W=8.8e-07 $X=71090 $Y=-6260 $D=4
M1512 VDD 670 Q2 VDD PM L=1.8e-07 W=8.8e-07 $X=71380 $Y=-19210 $D=4
M1513 VDD 671 Q7 VDD PM L=1.8e-07 W=8.8e-07 $X=71380 $Y=-3460 $D=4
M1514 277 673 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=72960 $Y=-42310 $D=4
M1515 276 674 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=72960 $Y=20080 $D=4
M1516 683 680 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=72990 $Y=-16410 $D=4
M1517 684 675 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=73030 $Y=-6260 $D=4
M1518 20 258 683 VDD PM L=1.8e-07 W=4.4e-07 $X=73750 $Y=-16410 $D=4
M1519 20 260 684 VDD PM L=1.8e-07 W=4.4e-07 $X=73790 $Y=-5820 $D=4
M1520 701 34 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=74080 $Y=-18770 $D=4
M1521 702 18 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=74080 $Y=-3460 $D=4
M1522 700 274 258 VDD PM L=1.8e-07 W=4.4e-07 $X=75840 $Y=-5820 $D=4
M1523 699 273 258 VDD PM L=1.8e-07 W=4.4e-07 $X=75890 $Y=-16410 $D=4
M1524 1503 CLK 695 VDD PM L=1.8e-07 W=8.8e-07 $X=76020 $Y=-19210 $D=4
M1525 1504 CLK 696 VDD PM L=1.8e-07 W=8.8e-07 $X=76020 $Y=-3460 $D=4
M1526 1505 RST 1503 VDD PM L=1.8e-07 W=8.8e-07 $X=76450 $Y=-19210 $D=4
M1527 1506 RST 1504 VDD PM L=1.8e-07 W=8.8e-07 $X=76450 $Y=-3460 $D=4
M1528 VDD 701 1505 VDD PM L=1.8e-07 W=8.8e-07 $X=76880 $Y=-19210 $D=4
M1529 VDD 702 1506 VDD PM L=1.8e-07 W=8.8e-07 $X=76880 $Y=-3460 $D=4
M1530 706 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=77600 $Y=-19210 $D=4
M1531 707 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=77600 $Y=-3460 $D=4
M1532 704 274 260 VDD PM L=1.8e-07 W=4.4e-07 $X=77790 $Y=-5820 $D=4
M1533 705 273 260 VDD PM L=1.8e-07 W=4.4e-07 $X=77830 $Y=-16410 $D=4
M1534 VDD 700 704 VDD PM L=1.8e-07 W=8.8e-07 $X=78550 $Y=-6260 $D=4
M1535 VDD 699 705 VDD PM L=1.8e-07 W=8.8e-07 $X=78590 $Y=-16410 $D=4
M1536 1507 272 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=79310 $Y=-16410 $D=4
M1537 700 263 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=79310 $Y=-5820 $D=4
M1538 699 263 1507 VDD PM L=1.8e-07 W=8.8e-07 $X=79740 $Y=-16410 $D=4
M1539 VDD 272 700 VDD PM L=1.8e-07 W=4.4e-07 $X=80030 $Y=-5820 $D=4
M1540 VDD 706 Q1 VDD PM L=1.8e-07 W=8.8e-07 $X=80300 $Y=-19210 $D=4
M1541 VDD 707 Q6 VDD PM L=1.8e-07 W=8.8e-07 $X=80300 $Y=-3460 $D=4
M1542 VDD 272 721 VDD PM L=1.8e-07 W=8.8e-07 $X=81680 $Y=-16410 $D=4
M1543 720 700 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=81970 $Y=-5820 $D=4
M1544 721 263 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=82400 $Y=-16410 $D=4
M1545 1508 263 720 VDD PM L=1.8e-07 W=8.8e-07 $X=82730 $Y=-6260 $D=4
M1546 748 35 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=83000 $Y=-18770 $D=4
M1547 749 29 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=83000 $Y=-3460 $D=4
M1548 732 699 721 VDD PM L=1.8e-07 W=8.8e-07 $X=83120 $Y=-16410 $D=4
M1549 VDD 272 1508 VDD PM L=1.8e-07 W=8.8e-07 $X=83160 $Y=-6260 $D=4
M1550 1509 CLK 734 VDD PM L=1.8e-07 W=8.8e-07 $X=84940 $Y=-19210 $D=4
M1551 1510 CLK 735 VDD PM L=1.8e-07 W=8.8e-07 $X=84940 $Y=-3460 $D=4
M1552 745 732 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=85060 $Y=-16410 $D=4
M1553 746 720 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=85100 $Y=-6260 $D=4
M1554 1511 RST 1509 VDD PM L=1.8e-07 W=8.8e-07 $X=85370 $Y=-19210 $D=4
M1555 1512 RST 1510 VDD PM L=1.8e-07 W=8.8e-07 $X=85370 $Y=-3460 $D=4
M1556 VDD 748 1511 VDD PM L=1.8e-07 W=8.8e-07 $X=85800 $Y=-19210 $D=4
M1557 VDD 749 1512 VDD PM L=1.8e-07 W=8.8e-07 $X=85800 $Y=-3460 $D=4
M1558 30 273 745 VDD PM L=1.8e-07 W=4.4e-07 $X=85820 $Y=-16410 $D=4
M1559 30 274 746 VDD PM L=1.8e-07 W=4.4e-07 $X=85860 $Y=-5820 $D=4
M1560 760 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=86520 $Y=-19210 $D=4
M1561 761 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=86520 $Y=-3460 $D=4
M1562 763 774 273 VDD PM L=1.8e-07 W=4.4e-07 $X=87910 $Y=-5820 $D=4
M1563 762 772 273 VDD PM L=1.8e-07 W=4.4e-07 $X=87960 $Y=-16410 $D=4
M1564 VDD 760 Q0 VDD PM L=1.8e-07 W=8.8e-07 $X=89220 $Y=-19210 $D=4
M1565 VDD 761 Q5 VDD PM L=1.8e-07 W=8.8e-07 $X=89220 $Y=-3460 $D=4
M1566 776 774 274 VDD PM L=1.8e-07 W=4.4e-07 $X=89860 $Y=-5820 $D=4
M1567 777 772 274 VDD PM L=1.8e-07 W=4.4e-07 $X=89900 $Y=-16410 $D=4
M1568 VDD 763 776 VDD PM L=1.8e-07 W=8.8e-07 $X=90620 $Y=-6260 $D=4
M1569 VDD 762 777 VDD PM L=1.8e-07 W=8.8e-07 $X=90660 $Y=-16410 $D=4
M1570 1513 277 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=91380 $Y=-16410 $D=4
M1571 763 276 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=91380 $Y=-5820 $D=4
M1572 762 276 1513 VDD PM L=1.8e-07 W=8.8e-07 $X=91810 $Y=-16410 $D=4
M1573 807 32 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=91920 $Y=-3460 $D=4
M1574 VDD 277 763 VDD PM L=1.8e-07 W=4.4e-07 $X=92100 $Y=-5820 $D=4
M1575 VDD 277 808 VDD PM L=1.8e-07 W=8.8e-07 $X=93750 $Y=-16410 $D=4
M1576 1514 CLK 789 VDD PM L=1.8e-07 W=8.8e-07 $X=93860 $Y=-3460 $D=4
M1577 806 763 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=94040 $Y=-5820 $D=4
M1578 1515 RST 1514 VDD PM L=1.8e-07 W=8.8e-07 $X=94290 $Y=-3460 $D=4
M1579 808 276 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=94470 $Y=-16410 $D=4
M1580 VDD 807 1515 VDD PM L=1.8e-07 W=8.8e-07 $X=94720 $Y=-3460 $D=4
M1581 1516 276 806 VDD PM L=1.8e-07 W=8.8e-07 $X=94800 $Y=-6260 $D=4
M1582 811 762 808 VDD PM L=1.8e-07 W=8.8e-07 $X=95190 $Y=-16410 $D=4
M1583 VDD 277 1516 VDD PM L=1.8e-07 W=8.8e-07 $X=95230 $Y=-6260 $D=4
M1584 813 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=95440 $Y=-3460 $D=4
M1585 VDD 264 817 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-135865 $D=4
M1586 VDD 265 818 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-133505 $D=4
M1587 VDD 266 819 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-120625 $D=4
M1588 VDD 267 820 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-118265 $D=4
M1589 VDD 268 821 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-105385 $D=4
M1590 VDD 269 822 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-103025 $D=4
M1591 VDD 270 823 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-90145 $D=4
M1592 VDD 271 824 VDD PM L=1.8e-07 W=8.8e-07 $X=96730 $Y=-87785 $D=4
M1593 815 811 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=97130 $Y=-16410 $D=4
M1594 816 806 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=97170 $Y=-6260 $D=4
M1595 34 772 815 VDD PM L=1.8e-07 W=4.4e-07 $X=97890 $Y=-16410 $D=4
M1596 34 774 816 VDD PM L=1.8e-07 W=4.4e-07 $X=97930 $Y=-5820 $D=4
M1597 VDD 813 Q4 VDD PM L=1.8e-07 W=8.8e-07 $X=98140 $Y=-3460 $D=4
M1598 VDD 826 836 VDD PM L=1.8e-07 W=8.8e-07 $X=99510 $Y=-74905 $D=4
M1599 VDD 772 774 VDD PM L=1.8e-07 W=4.4e-07 $X=99950 $Y=-5820 $D=4
M1600 772 278 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=100670 $Y=-5820 $D=4
M1601 VDD 828 838 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-135865 $D=4
M1602 VDD 829 839 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-133505 $D=4
M1603 VDD 830 840 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-120625 $D=4
M1604 VDD 831 841 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-118265 $D=4
M1605 VDD 832 842 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-105385 $D=4
M1606 VDD 833 843 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-103025 $D=4
M1607 VDD 834 844 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-90145 $D=4
M1608 VDD 835 845 VDD PM L=1.8e-07 W=8.8e-07 $X=101370 $Y=-87785 $D=4
M1609 VDD 283 772 VDD PM L=1.8e-07 W=4.4e-07 $X=101390 $Y=-5820 $D=4
M1610 837 827 VDD VDD PM L=1.8e-07 W=1.76e-06 $X=102250 $Y=-151985 $D=4
M1611 846 772 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=103330 $Y=-5820 $D=4
M1612 281 GND VDD VDD PM L=1.8e-07 W=4.4e-07 $X=103470 $Y=-148745 $D=4
M1613 1517 278 846 VDD PM L=1.8e-07 W=8.8e-07 $X=104090 $Y=-6260 $D=4
M1614 VDD 283 1517 VDD PM L=1.8e-07 W=8.8e-07 $X=104520 $Y=-6260 $D=4
M1615 857 856 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=106170 $Y=-150665 $D=4
M1616 35 846 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=106460 $Y=-5820 $D=4
M1617 261 279 1518 VDD PM L=1.8e-07 W=8.8e-07 $X=107900 $Y=-148745 $D=4
M1618 1519 281 261 VDD PM L=1.8e-07 W=8.8e-07 $X=108620 $Y=-148745 $D=4
M1619 1520 282 262 VDD PM L=1.8e-07 W=8.8e-07 $X=108620 $Y=-74905 $D=4
M1620 VDD 857 858 VDD PM L=1.8e-07 W=8.8e-07 $X=108870 $Y=-151105 $D=4
M1621 VDD 292 1519 VDD PM L=1.8e-07 W=8.8e-07 $X=109050 $Y=-148745 $D=4
M1622 VDD 293 1520 VDD PM L=1.8e-07 W=8.8e-07 $X=109050 $Y=-74905 $D=4
M1623 1521 294 866 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-135865 $D=4
M1624 1522 295 867 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-133505 $D=4
M1625 1523 296 868 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-120625 $D=4
M1626 1524 297 863 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-118265 $D=4
M1627 1525 298 864 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-105385 $D=4
M1628 1526 299 869 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-103025 $D=4
M1629 1527 300 870 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-90145 $D=4
M1630 1528 301 871 VDD PM L=1.8e-07 W=8.8e-07 $X=112500 $Y=-87785 $D=4
M1631 VDD 305 1521 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-135865 $D=4
M1632 VDD 306 1522 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-133505 $D=4
M1633 VDD 307 1523 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-120625 $D=4
M1634 VDD 308 1524 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-118265 $D=4
M1635 VDD 309 1525 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-105385 $D=4
M1636 VDD 310 1526 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-103025 $D=4
M1637 VDD 311 1527 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-90145 $D=4
M1638 VDD 312 1528 VDD PM L=1.8e-07 W=8.8e-07 $X=112930 $Y=-87785 $D=4
M1639 7 894 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=118450 $Y=-168225 $D=4
M1640 8 895 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=118450 $Y=-158075 $D=4
M1641 VDD 37 322 VDD PM L=1.8e-07 W=4.4e-07 $X=119100 $Y=-146485 $D=4
M1642 VDD 874 874 VDD PM L=1.8e-07 W=3.3e-06 $X=119100 $Y=-137205 $D=4
M1643 326 322 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=119820 $Y=-146485 $D=4
M1644 VDD 323 894 VDD PM L=1.8e-07 W=8.8e-07 $X=121150 $Y=-168225 $D=4
M1645 VDD 323 895 VDD PM L=1.8e-07 W=8.8e-07 $X=121150 $Y=-158075 $D=4
M1646 1529 910 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=121870 $Y=-168225 $D=4
M1647 1530 911 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=121870 $Y=-158075 $D=4
M1648 1531 RST 1529 VDD PM L=1.8e-07 W=8.8e-07 $X=122300 $Y=-168225 $D=4
M1649 1532 RST 1530 VDD PM L=1.8e-07 W=8.8e-07 $X=122300 $Y=-158075 $D=4
M1650 898 323 1531 VDD PM L=1.8e-07 W=8.8e-07 $X=122730 $Y=-168225 $D=4
M1651 899 323 1532 VDD PM L=1.8e-07 W=8.8e-07 $X=122730 $Y=-158075 $D=4
M1652 VDD 38 327 VDD PM L=1.8e-07 W=4.4e-07 $X=123560 $Y=-146485 $D=4
M1653 VDD 900 900 VDD PM L=1.8e-07 W=3.3e-06 $X=123560 $Y=-137205 $D=4
M1654 330 327 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=124280 $Y=-146485 $D=4
M1655 VDD 39 910 VDD PM L=1.8e-07 W=4.4e-07 $X=124670 $Y=-168225 $D=4
M1656 VDD 36 911 VDD PM L=1.8e-07 W=4.4e-07 $X=124670 $Y=-157635 $D=4
M1657 11 934 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=126650 $Y=-168225 $D=4
M1658 9 935 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=126650 $Y=-158075 $D=4
M1659 VDD 41 331 VDD PM L=1.8e-07 W=4.4e-07 $X=128020 $Y=-146485 $D=4
M1660 VDD 924 924 VDD PM L=1.8e-07 W=3.3e-06 $X=128020 $Y=-137205 $D=4
M1661 334 331 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=128740 $Y=-146485 $D=4
M1662 VDD 323 934 VDD PM L=1.8e-07 W=8.8e-07 $X=129350 $Y=-168225 $D=4
M1663 VDD 323 935 VDD PM L=1.8e-07 W=8.8e-07 $X=129350 $Y=-158075 $D=4
M1664 1533 959 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=130070 $Y=-168225 $D=4
M1665 1534 960 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=130070 $Y=-158075 $D=4
M1666 1535 RST 1533 VDD PM L=1.8e-07 W=8.8e-07 $X=130500 $Y=-168225 $D=4
M1667 1536 RST 1534 VDD PM L=1.8e-07 W=8.8e-07 $X=130500 $Y=-158075 $D=4
M1668 948 323 1535 VDD PM L=1.8e-07 W=8.8e-07 $X=130930 $Y=-168225 $D=4
M1669 949 323 1536 VDD PM L=1.8e-07 W=8.8e-07 $X=130930 $Y=-158075 $D=4
M1670 VDD 42 335 VDD PM L=1.8e-07 W=4.4e-07 $X=132480 $Y=-146485 $D=4
M1671 VDD 950 950 VDD PM L=1.8e-07 W=3.3e-06 $X=132480 $Y=-137205 $D=4
M1672 VDD 43 959 VDD PM L=1.8e-07 W=4.4e-07 $X=132870 $Y=-168225 $D=4
M1673 VDD 40 960 VDD PM L=1.8e-07 W=4.4e-07 $X=132870 $Y=-157635 $D=4
M1674 338 335 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=133200 $Y=-146485 $D=4
M1675 12 983 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=134850 $Y=-168225 $D=4
M1676 13 984 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=134850 $Y=-158075 $D=4
M1677 VDD 45 339 VDD PM L=1.8e-07 W=4.4e-07 $X=136940 $Y=-146485 $D=4
M1678 VDD 974 974 VDD PM L=1.8e-07 W=3.3e-06 $X=136940 $Y=-137205 $D=4
M1679 VDD 323 983 VDD PM L=1.8e-07 W=8.8e-07 $X=137550 $Y=-168225 $D=4
M1680 VDD 323 984 VDD PM L=1.8e-07 W=8.8e-07 $X=137550 $Y=-158075 $D=4
M1681 342 339 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=137660 $Y=-146485 $D=4
M1682 1537 1000 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=138270 $Y=-168225 $D=4
M1683 1538 1001 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=138270 $Y=-158075 $D=4
M1684 1539 RST 1537 VDD PM L=1.8e-07 W=8.8e-07 $X=138700 $Y=-168225 $D=4
M1685 1540 RST 1538 VDD PM L=1.8e-07 W=8.8e-07 $X=138700 $Y=-158075 $D=4
M1686 997 323 1539 VDD PM L=1.8e-07 W=8.8e-07 $X=139130 $Y=-168225 $D=4
M1687 998 323 1540 VDD PM L=1.8e-07 W=8.8e-07 $X=139130 $Y=-158075 $D=4
M1688 VDD 46 1000 VDD PM L=1.8e-07 W=4.4e-07 $X=141070 $Y=-168225 $D=4
M1689 VDD 44 1001 VDD PM L=1.8e-07 W=4.4e-07 $X=141070 $Y=-157635 $D=4
M1690 VDD 47 343 VDD PM L=1.8e-07 W=4.4e-07 $X=141400 $Y=-146485 $D=4
M1691 VDD 1002 1002 VDD PM L=1.8e-07 W=3.3e-06 $X=141400 $Y=-137205 $D=4
M1692 346 343 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=142120 $Y=-146485 $D=4
M1693 6 1024 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=143050 $Y=-168225 $D=4
M1694 10 1025 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=143050 $Y=-158075 $D=4
M1695 VDD 323 1024 VDD PM L=1.8e-07 W=8.8e-07 $X=145750 $Y=-168225 $D=4
M1696 VDD 323 1025 VDD PM L=1.8e-07 W=8.8e-07 $X=145750 $Y=-158075 $D=4
M1697 VDD 49 347 VDD PM L=1.8e-07 W=4.4e-07 $X=145860 $Y=-146485 $D=4
M1698 VDD 1026 1026 VDD PM L=1.8e-07 W=3.3e-06 $X=145860 $Y=-137205 $D=4
M1699 1541 1049 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=146470 $Y=-168225 $D=4
M1700 1542 1050 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=146470 $Y=-158075 $D=4
M1701 350 347 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=146580 $Y=-146485 $D=4
M1702 1543 RST 1541 VDD PM L=1.8e-07 W=8.8e-07 $X=146900 $Y=-168225 $D=4
M1703 1544 RST 1542 VDD PM L=1.8e-07 W=8.8e-07 $X=146900 $Y=-158075 $D=4
M1704 1047 323 1543 VDD PM L=1.8e-07 W=8.8e-07 $X=147330 $Y=-168225 $D=4
M1705 1048 323 1544 VDD PM L=1.8e-07 W=8.8e-07 $X=147330 $Y=-158075 $D=4
M1706 VDD 51 1049 VDD PM L=1.8e-07 W=4.4e-07 $X=149270 $Y=-168225 $D=4
M1707 VDD 48 1050 VDD PM L=1.8e-07 W=4.4e-07 $X=149270 $Y=-157635 $D=4
M1708 VDD 52 351 VDD PM L=1.8e-07 W=4.4e-07 $X=150320 $Y=-146485 $D=4
M1709 VDD 1052 1052 VDD PM L=1.8e-07 W=3.3e-06 $X=150320 $Y=-137205 $D=4
M1710 354 351 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=151040 $Y=-146485 $D=4
M1711 53 1073 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=151250 $Y=-168225 $D=4
M1712 54 1074 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=151250 $Y=-158075 $D=4
M1713 VDD 323 1073 VDD PM L=1.8e-07 W=8.8e-07 $X=153950 $Y=-168225 $D=4
M1714 VDD 323 1074 VDD PM L=1.8e-07 W=8.8e-07 $X=153950 $Y=-158075 $D=4
M1715 1545 1099 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=154670 $Y=-168225 $D=4
M1716 1546 1100 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=154670 $Y=-158075 $D=4
M1717 VDD 56 355 VDD PM L=1.8e-07 W=4.4e-07 $X=154780 $Y=-146485 $D=4
M1718 VDD 1076 1076 VDD PM L=1.8e-07 W=3.3e-06 $X=154780 $Y=-137205 $D=4
M1719 1547 RST 1545 VDD PM L=1.8e-07 W=8.8e-07 $X=155100 $Y=-168225 $D=4
M1720 1548 RST 1546 VDD PM L=1.8e-07 W=8.8e-07 $X=155100 $Y=-158075 $D=4
M1721 358 355 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=155500 $Y=-146485 $D=4
M1722 1095 323 1547 VDD PM L=1.8e-07 W=8.8e-07 $X=155530 $Y=-168225 $D=4
M1723 1096 323 1548 VDD PM L=1.8e-07 W=8.8e-07 $X=155530 $Y=-158075 $D=4
M1724 VDD 57 1099 VDD PM L=1.8e-07 W=4.4e-07 $X=157470 $Y=-168225 $D=4
M1725 VDD 55 1100 VDD PM L=1.8e-07 W=4.4e-07 $X=157470 $Y=-157635 $D=4
M1726 VDD 58 359 VDD PM L=1.8e-07 W=4.4e-07 $X=159240 $Y=-146485 $D=4
M1727 VDD 1102 1102 VDD PM L=1.8e-07 W=3.3e-06 $X=159240 $Y=-137205 $D=4
M1728 59 1123 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=159450 $Y=-168225 $D=4
M1729 61 1124 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=159450 $Y=-158075 $D=4
M1730 362 359 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=159960 $Y=-146485 $D=4
M1731 VDD 323 1123 VDD PM L=1.8e-07 W=8.8e-07 $X=162150 $Y=-168225 $D=4
M1732 VDD 323 1124 VDD PM L=1.8e-07 W=8.8e-07 $X=162150 $Y=-158075 $D=4
M1733 1549 1148 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=162870 $Y=-168225 $D=4
M1734 1550 1149 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=162870 $Y=-158075 $D=4
M1735 1551 RST 1549 VDD PM L=1.8e-07 W=8.8e-07 $X=163300 $Y=-168225 $D=4
M1736 1552 RST 1550 VDD PM L=1.8e-07 W=8.8e-07 $X=163300 $Y=-158075 $D=4
M1737 VDD 62 363 VDD PM L=1.8e-07 W=4.4e-07 $X=163700 $Y=-146485 $D=4
M1738 VDD 1126 1126 VDD PM L=1.8e-07 W=3.3e-06 $X=163700 $Y=-137205 $D=4
M1739 1136 323 1551 VDD PM L=1.8e-07 W=8.8e-07 $X=163730 $Y=-168225 $D=4
M1740 1137 323 1552 VDD PM L=1.8e-07 W=8.8e-07 $X=163730 $Y=-158075 $D=4
M1741 366 363 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=164420 $Y=-146485 $D=4
M1742 VDD 64 1148 VDD PM L=1.8e-07 W=4.4e-07 $X=165670 $Y=-168225 $D=4
M1743 VDD 60 1149 VDD PM L=1.8e-07 W=4.4e-07 $X=165670 $Y=-157635 $D=4
M1744 63 1173 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=167650 $Y=-168225 $D=4
M1745 65 1174 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=167650 $Y=-158075 $D=4
M1746 VDD 66 367 VDD PM L=1.8e-07 W=4.4e-07 $X=168160 $Y=-146485 $D=4
M1747 VDD 1152 1152 VDD PM L=1.8e-07 W=3.3e-06 $X=168160 $Y=-137205 $D=4
M1748 370 367 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=168880 $Y=-146485 $D=4
M1749 VDD 323 1173 VDD PM L=1.8e-07 W=8.8e-07 $X=170350 $Y=-168225 $D=4
M1750 VDD 323 1174 VDD PM L=1.8e-07 W=8.8e-07 $X=170350 $Y=-158075 $D=4
M1751 1553 1188 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=171070 $Y=-168225 $D=4
M1752 1554 1189 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=171070 $Y=-158075 $D=4
M1753 1555 RST 1553 VDD PM L=1.8e-07 W=8.8e-07 $X=171500 $Y=-168225 $D=4
M1754 1556 RST 1554 VDD PM L=1.8e-07 W=8.8e-07 $X=171500 $Y=-158075 $D=4
M1755 1177 323 1555 VDD PM L=1.8e-07 W=8.8e-07 $X=171930 $Y=-168225 $D=4
M1756 1178 323 1556 VDD PM L=1.8e-07 W=8.8e-07 $X=171930 $Y=-158075 $D=4
M1757 VDD 68 371 VDD PM L=1.8e-07 W=4.4e-07 $X=172620 $Y=-146485 $D=4
M1758 VDD 1176 1176 VDD PM L=1.8e-07 W=3.3e-06 $X=172620 $Y=-137205 $D=4
M1759 374 371 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=173340 $Y=-146485 $D=4
M1760 VDD 69 1188 VDD PM L=1.8e-07 W=4.4e-07 $X=173870 $Y=-168225 $D=4
M1761 VDD 67 1189 VDD PM L=1.8e-07 W=4.4e-07 $X=173870 $Y=-157635 $D=4
M1762 70 1221 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=175850 $Y=-168225 $D=4
M1763 73 1222 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=175850 $Y=-158075 $D=4
M1764 VDD 71 375 VDD PM L=1.8e-07 W=4.4e-07 $X=177080 $Y=-146485 $D=4
M1765 VDD 1202 1202 VDD PM L=1.8e-07 W=3.3e-06 $X=177080 $Y=-137205 $D=4
M1766 378 375 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=177800 $Y=-146485 $D=4
M1767 VDD 323 1221 VDD PM L=1.8e-07 W=8.8e-07 $X=178550 $Y=-168225 $D=4
M1768 VDD 323 1222 VDD PM L=1.8e-07 W=8.8e-07 $X=178550 $Y=-158075 $D=4
M1769 1557 1237 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=179270 $Y=-168225 $D=4
M1770 1558 1238 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=179270 $Y=-158075 $D=4
M1771 1559 RST 1557 VDD PM L=1.8e-07 W=8.8e-07 $X=179700 $Y=-168225 $D=4
M1772 1560 RST 1558 VDD PM L=1.8e-07 W=8.8e-07 $X=179700 $Y=-158075 $D=4
M1773 1226 323 1559 VDD PM L=1.8e-07 W=8.8e-07 $X=180130 $Y=-168225 $D=4
M1774 1227 323 1560 VDD PM L=1.8e-07 W=8.8e-07 $X=180130 $Y=-158075 $D=4
M1775 VDD 74 379 VDD PM L=1.8e-07 W=4.4e-07 $X=181540 $Y=-146485 $D=4
M1776 VDD 1228 1228 VDD PM L=1.8e-07 W=3.3e-06 $X=181540 $Y=-137205 $D=4
M1777 VDD 75 1237 VDD PM L=1.8e-07 W=4.4e-07 $X=182070 $Y=-168225 $D=4
M1778 VDD 72 1238 VDD PM L=1.8e-07 W=4.4e-07 $X=182070 $Y=-157635 $D=4
M1779 382 379 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=182260 $Y=-146485 $D=4
M1780 VDD 76 383 VDD PM L=1.8e-07 W=4.4e-07 $X=186000 $Y=-146485 $D=4
M1781 VDD 1252 1252 VDD PM L=1.8e-07 W=3.3e-06 $X=186000 $Y=-137205 $D=4
M1782 386 383 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=186720 $Y=-146485 $D=4
X1783 GND 893 883 325 n18_CDNS_6738901947925 $T=120000 -139615 1 180 $X=119160 $Y=-139965
X1784 GND 921 909 329 n18_CDNS_6738901947925 $T=124460 -139615 1 180 $X=123620 $Y=-139965
X1785 GND 945 933 333 n18_CDNS_6738901947925 $T=128920 -139615 1 180 $X=128080 $Y=-139965
X1786 GND 971 961 337 n18_CDNS_6738901947925 $T=133380 -139615 1 180 $X=132540 $Y=-139965
X1787 GND 995 985 341 n18_CDNS_6738901947925 $T=137840 -139615 1 180 $X=137000 $Y=-139965
X1788 GND 1021 1011 345 n18_CDNS_6738901947925 $T=142300 -139615 1 180 $X=141460 $Y=-139965
X1789 GND 1045 1035 349 n18_CDNS_6738901947925 $T=146760 -139615 1 180 $X=145920 $Y=-139965
X1790 GND 1071 1061 353 n18_CDNS_6738901947925 $T=151220 -139615 1 180 $X=150380 $Y=-139965
X1791 GND 1097 1085 357 n18_CDNS_6738901947925 $T=155680 -139615 1 180 $X=154840 $Y=-139965
X1792 GND 1121 1111 361 n18_CDNS_6738901947925 $T=160140 -139615 1 180 $X=159300 $Y=-139965
X1793 GND 1147 1135 365 n18_CDNS_6738901947925 $T=164600 -139615 1 180 $X=163760 $Y=-139965
X1794 GND 1171 1161 369 n18_CDNS_6738901947925 $T=169060 -139615 1 180 $X=168220 $Y=-139965
X1795 GND 1199 1187 373 n18_CDNS_6738901947925 $T=173520 -139615 1 180 $X=172680 $Y=-139965
X1796 GND 1223 1211 377 n18_CDNS_6738901947925 $T=177980 -139615 1 180 $X=177140 $Y=-139965
X1797 GND 1249 1239 381 n18_CDNS_6738901947925 $T=182440 -139615 1 180 $X=181600 $Y=-139965
X1798 GND 1271 1261 385 n18_CDNS_6738901947925 $T=186900 -139615 1 180 $X=186060 $Y=-139965
X1799 VDD 893 874 p18_CDNS_6738901947922 $T=120000 -137205 1 180 $X=118910 $Y=-137635
X1800 VDD 921 900 p18_CDNS_6738901947922 $T=124460 -137205 1 180 $X=123370 $Y=-137635
X1801 VDD 945 924 p18_CDNS_6738901947922 $T=128920 -137205 1 180 $X=127830 $Y=-137635
X1802 VDD 971 950 p18_CDNS_6738901947922 $T=133380 -137205 1 180 $X=132290 $Y=-137635
X1803 VDD 995 974 p18_CDNS_6738901947922 $T=137840 -137205 1 180 $X=136750 $Y=-137635
X1804 VDD 1021 1002 p18_CDNS_6738901947922 $T=142300 -137205 1 180 $X=141210 $Y=-137635
X1805 VDD 1045 1026 p18_CDNS_6738901947922 $T=146760 -137205 1 180 $X=145670 $Y=-137635
X1806 VDD 1071 1052 p18_CDNS_6738901947922 $T=151220 -137205 1 180 $X=150130 $Y=-137635
X1807 VDD 1097 1076 p18_CDNS_6738901947922 $T=155680 -137205 1 180 $X=154590 $Y=-137635
X1808 VDD 1121 1102 p18_CDNS_6738901947922 $T=160140 -137205 1 180 $X=159050 $Y=-137635
X1809 VDD 1147 1126 p18_CDNS_6738901947922 $T=164600 -137205 1 180 $X=163510 $Y=-137635
X1810 VDD 1171 1152 p18_CDNS_6738901947922 $T=169060 -137205 1 180 $X=167970 $Y=-137635
X1811 VDD 1199 1176 p18_CDNS_6738901947922 $T=173520 -137205 1 180 $X=172430 $Y=-137635
X1812 VDD 1223 1202 p18_CDNS_6738901947922 $T=177980 -137205 1 180 $X=176890 $Y=-137635
X1813 VDD 1249 1228 p18_CDNS_6738901947922 $T=182440 -137205 1 180 $X=181350 $Y=-137635
X1814 VDD 1271 1252 p18_CDNS_6738901947922 $T=186900 -137205 1 180 $X=185810 $Y=-137635
X1815 324 325 873 VDD p18_CDNS_6738901947929 $T=119330 -83535 0 270 $X=118900 $Y=-84625
X1816 328 329 873 VDD p18_CDNS_6738901947929 $T=123790 -83535 0 270 $X=123360 $Y=-84625
X1817 332 333 873 VDD p18_CDNS_6738901947929 $T=128250 -83535 0 270 $X=127820 $Y=-84625
X1818 336 337 873 VDD p18_CDNS_6738901947929 $T=132710 -83535 0 270 $X=132280 $Y=-84625
X1819 340 341 873 VDD p18_CDNS_6738901947929 $T=137170 -83535 0 270 $X=136740 $Y=-84625
X1820 344 345 873 VDD p18_CDNS_6738901947929 $T=141630 -83535 0 270 $X=141200 $Y=-84625
X1821 348 349 873 VDD p18_CDNS_6738901947929 $T=146090 -83535 0 270 $X=145660 $Y=-84625
X1822 352 353 873 VDD p18_CDNS_6738901947929 $T=150550 -83535 0 270 $X=150120 $Y=-84625
X1823 356 357 873 VDD p18_CDNS_6738901947929 $T=155010 -83535 0 270 $X=154580 $Y=-84625
X1824 360 361 873 VDD p18_CDNS_6738901947929 $T=159470 -83535 0 270 $X=159040 $Y=-84625
X1825 364 365 873 VDD p18_CDNS_6738901947929 $T=163930 -83535 0 270 $X=163500 $Y=-84625
X1826 368 369 873 VDD p18_CDNS_6738901947929 $T=168390 -83535 0 270 $X=167960 $Y=-84625
X1827 372 373 873 VDD p18_CDNS_6738901947929 $T=172850 -83535 0 270 $X=172420 $Y=-84625
X1828 376 377 873 VDD p18_CDNS_6738901947929 $T=177310 -83535 0 270 $X=176880 $Y=-84625
X1829 380 381 873 VDD p18_CDNS_6738901947929 $T=181770 -83535 0 270 $X=181340 $Y=-84625
X1830 384 385 873 VDD p18_CDNS_6738901947929 $T=186230 -83535 0 270 $X=185800 $Y=-84625
X1831 GND 883 865 n18_CDNS_6738901947921 $T=119110 -141245 1 90 $X=118760 $Y=-141905
X1832 GND 909 865 n18_CDNS_6738901947921 $T=123570 -141245 1 90 $X=123220 $Y=-141905
X1833 GND 933 865 n18_CDNS_6738901947921 $T=128030 -141245 1 90 $X=127680 $Y=-141905
X1834 GND 961 865 n18_CDNS_6738901947921 $T=132490 -141245 1 90 $X=132140 $Y=-141905
X1835 GND 985 865 n18_CDNS_6738901947921 $T=136950 -141245 1 90 $X=136600 $Y=-141905
X1836 GND 1011 865 n18_CDNS_6738901947921 $T=141410 -141245 1 90 $X=141060 $Y=-141905
X1837 GND 1035 865 n18_CDNS_6738901947921 $T=145870 -141245 1 90 $X=145520 $Y=-141905
X1838 GND 1061 865 n18_CDNS_6738901947921 $T=150330 -141245 1 90 $X=149980 $Y=-141905
X1839 GND 1085 865 n18_CDNS_6738901947921 $T=154790 -141245 1 90 $X=154440 $Y=-141905
X1840 GND 1111 865 n18_CDNS_6738901947921 $T=159250 -141245 1 90 $X=158900 $Y=-141905
X1841 GND 1135 865 n18_CDNS_6738901947921 $T=163710 -141245 1 90 $X=163360 $Y=-141905
X1842 GND 1161 865 n18_CDNS_6738901947921 $T=168170 -141245 1 90 $X=167820 $Y=-141905
X1843 GND 1187 865 n18_CDNS_6738901947921 $T=172630 -141245 1 90 $X=172280 $Y=-141905
X1844 GND 1211 865 n18_CDNS_6738901947921 $T=177090 -141245 1 90 $X=176740 $Y=-141905
X1845 GND 1239 865 n18_CDNS_6738901947921 $T=181550 -141245 1 90 $X=181200 $Y=-141905
X1846 GND 1261 865 n18_CDNS_6738901947921 $T=186010 -141245 1 90 $X=185660 $Y=-141905
X1847 325 885 324 875 866 GND ICV_1 $T=118940 -131675 0 90 $X=118150 $Y=-132335
X1848 325 886 324 876 867 GND ICV_1 $T=118940 -125635 0 90 $X=118150 $Y=-126295
X1849 325 887 324 877 868 GND ICV_1 $T=118940 -119595 0 90 $X=118150 $Y=-120255
X1850 325 888 324 878 863 GND ICV_1 $T=118940 -113555 0 90 $X=118150 $Y=-114215
X1851 325 889 324 879 864 GND ICV_1 $T=118940 -107515 0 90 $X=118150 $Y=-108175
X1852 325 890 324 880 869 GND ICV_1 $T=118940 -101475 0 90 $X=118150 $Y=-102135
X1853 325 891 324 881 870 GND ICV_1 $T=118940 -95435 0 90 $X=118150 $Y=-96095
X1854 325 892 324 882 871 GND ICV_1 $T=118940 -89395 0 90 $X=118150 $Y=-90055
X1855 329 913 328 901 866 GND ICV_1 $T=123400 -131675 0 90 $X=122610 $Y=-132335
X1856 329 914 328 902 867 GND ICV_1 $T=123400 -125635 0 90 $X=122610 $Y=-126295
X1857 329 915 328 903 868 GND ICV_1 $T=123400 -119595 0 90 $X=122610 $Y=-120255
X1858 329 916 328 904 863 GND ICV_1 $T=123400 -113555 0 90 $X=122610 $Y=-114215
X1859 329 917 328 905 864 GND ICV_1 $T=123400 -107515 0 90 $X=122610 $Y=-108175
X1860 329 918 328 906 869 GND ICV_1 $T=123400 -101475 0 90 $X=122610 $Y=-102135
X1861 329 919 328 907 870 GND ICV_1 $T=123400 -95435 0 90 $X=122610 $Y=-96095
X1862 329 920 328 908 871 GND ICV_1 $T=123400 -89395 0 90 $X=122610 $Y=-90055
X1863 333 937 332 925 866 GND ICV_1 $T=127860 -131675 0 90 $X=127070 $Y=-132335
X1864 333 938 332 926 867 GND ICV_1 $T=127860 -125635 0 90 $X=127070 $Y=-126295
X1865 333 939 332 927 868 GND ICV_1 $T=127860 -119595 0 90 $X=127070 $Y=-120255
X1866 333 940 332 928 863 GND ICV_1 $T=127860 -113555 0 90 $X=127070 $Y=-114215
X1867 333 941 332 929 864 GND ICV_1 $T=127860 -107515 0 90 $X=127070 $Y=-108175
X1868 333 942 332 930 869 GND ICV_1 $T=127860 -101475 0 90 $X=127070 $Y=-102135
X1869 333 943 332 931 870 GND ICV_1 $T=127860 -95435 0 90 $X=127070 $Y=-96095
X1870 333 944 332 932 871 GND ICV_1 $T=127860 -89395 0 90 $X=127070 $Y=-90055
X1871 337 963 336 951 866 GND ICV_1 $T=132320 -131675 0 90 $X=131530 $Y=-132335
X1872 337 964 336 952 867 GND ICV_1 $T=132320 -125635 0 90 $X=131530 $Y=-126295
X1873 337 965 336 953 868 GND ICV_1 $T=132320 -119595 0 90 $X=131530 $Y=-120255
X1874 337 966 336 954 863 GND ICV_1 $T=132320 -113555 0 90 $X=131530 $Y=-114215
X1875 337 967 336 955 864 GND ICV_1 $T=132320 -107515 0 90 $X=131530 $Y=-108175
X1876 337 968 336 956 869 GND ICV_1 $T=132320 -101475 0 90 $X=131530 $Y=-102135
X1877 337 969 336 957 870 GND ICV_1 $T=132320 -95435 0 90 $X=131530 $Y=-96095
X1878 337 970 336 958 871 GND ICV_1 $T=132320 -89395 0 90 $X=131530 $Y=-90055
X1879 341 987 340 975 866 GND ICV_1 $T=136780 -131675 0 90 $X=135990 $Y=-132335
X1880 341 988 340 976 867 GND ICV_1 $T=136780 -125635 0 90 $X=135990 $Y=-126295
X1881 341 989 340 977 868 GND ICV_1 $T=136780 -119595 0 90 $X=135990 $Y=-120255
X1882 341 990 340 978 863 GND ICV_1 $T=136780 -113555 0 90 $X=135990 $Y=-114215
X1883 341 991 340 979 864 GND ICV_1 $T=136780 -107515 0 90 $X=135990 $Y=-108175
X1884 341 992 340 980 869 GND ICV_1 $T=136780 -101475 0 90 $X=135990 $Y=-102135
X1885 341 993 340 981 870 GND ICV_1 $T=136780 -95435 0 90 $X=135990 $Y=-96095
X1886 341 994 340 982 871 GND ICV_1 $T=136780 -89395 0 90 $X=135990 $Y=-90055
X1887 345 1013 344 1003 866 GND ICV_1 $T=141240 -131675 0 90 $X=140450 $Y=-132335
X1888 345 1014 344 1004 867 GND ICV_1 $T=141240 -125635 0 90 $X=140450 $Y=-126295
X1889 345 1015 344 1005 868 GND ICV_1 $T=141240 -119595 0 90 $X=140450 $Y=-120255
X1890 345 1016 344 1006 863 GND ICV_1 $T=141240 -113555 0 90 $X=140450 $Y=-114215
X1891 345 1017 344 1007 864 GND ICV_1 $T=141240 -107515 0 90 $X=140450 $Y=-108175
X1892 345 1018 344 1008 869 GND ICV_1 $T=141240 -101475 0 90 $X=140450 $Y=-102135
X1893 345 1019 344 1009 870 GND ICV_1 $T=141240 -95435 0 90 $X=140450 $Y=-96095
X1894 345 1020 344 1010 871 GND ICV_1 $T=141240 -89395 0 90 $X=140450 $Y=-90055
X1895 349 1037 348 1027 866 GND ICV_1 $T=145700 -131675 0 90 $X=144910 $Y=-132335
X1896 349 1038 348 1028 867 GND ICV_1 $T=145700 -125635 0 90 $X=144910 $Y=-126295
X1897 349 1039 348 1029 868 GND ICV_1 $T=145700 -119595 0 90 $X=144910 $Y=-120255
X1898 349 1040 348 1030 863 GND ICV_1 $T=145700 -113555 0 90 $X=144910 $Y=-114215
X1899 349 1041 348 1031 864 GND ICV_1 $T=145700 -107515 0 90 $X=144910 $Y=-108175
X1900 349 1042 348 1032 869 GND ICV_1 $T=145700 -101475 0 90 $X=144910 $Y=-102135
X1901 349 1043 348 1033 870 GND ICV_1 $T=145700 -95435 0 90 $X=144910 $Y=-96095
X1902 349 1044 348 1034 871 GND ICV_1 $T=145700 -89395 0 90 $X=144910 $Y=-90055
X1903 353 1063 352 1053 866 GND ICV_1 $T=150160 -131675 0 90 $X=149370 $Y=-132335
X1904 353 1064 352 1054 867 GND ICV_1 $T=150160 -125635 0 90 $X=149370 $Y=-126295
X1905 353 1065 352 1055 868 GND ICV_1 $T=150160 -119595 0 90 $X=149370 $Y=-120255
X1906 353 1066 352 1056 863 GND ICV_1 $T=150160 -113555 0 90 $X=149370 $Y=-114215
X1907 353 1067 352 1057 864 GND ICV_1 $T=150160 -107515 0 90 $X=149370 $Y=-108175
X1908 353 1068 352 1058 869 GND ICV_1 $T=150160 -101475 0 90 $X=149370 $Y=-102135
X1909 353 1069 352 1059 870 GND ICV_1 $T=150160 -95435 0 90 $X=149370 $Y=-96095
X1910 353 1070 352 1060 871 GND ICV_1 $T=150160 -89395 0 90 $X=149370 $Y=-90055
X1911 357 1087 356 1077 866 GND ICV_1 $T=154620 -131675 0 90 $X=153830 $Y=-132335
X1912 357 1088 356 1078 867 GND ICV_1 $T=154620 -125635 0 90 $X=153830 $Y=-126295
X1913 357 1089 356 1079 868 GND ICV_1 $T=154620 -119595 0 90 $X=153830 $Y=-120255
X1914 357 1090 356 1080 863 GND ICV_1 $T=154620 -113555 0 90 $X=153830 $Y=-114215
X1915 357 1091 356 1081 864 GND ICV_1 $T=154620 -107515 0 90 $X=153830 $Y=-108175
X1916 357 1092 356 1082 869 GND ICV_1 $T=154620 -101475 0 90 $X=153830 $Y=-102135
X1917 357 1093 356 1083 870 GND ICV_1 $T=154620 -95435 0 90 $X=153830 $Y=-96095
X1918 357 1094 356 1084 871 GND ICV_1 $T=154620 -89395 0 90 $X=153830 $Y=-90055
X1919 361 1113 360 1103 866 GND ICV_1 $T=159080 -131675 0 90 $X=158290 $Y=-132335
X1920 361 1114 360 1104 867 GND ICV_1 $T=159080 -125635 0 90 $X=158290 $Y=-126295
X1921 361 1115 360 1105 868 GND ICV_1 $T=159080 -119595 0 90 $X=158290 $Y=-120255
X1922 361 1116 360 1106 863 GND ICV_1 $T=159080 -113555 0 90 $X=158290 $Y=-114215
X1923 361 1117 360 1107 864 GND ICV_1 $T=159080 -107515 0 90 $X=158290 $Y=-108175
X1924 361 1118 360 1108 869 GND ICV_1 $T=159080 -101475 0 90 $X=158290 $Y=-102135
X1925 361 1119 360 1109 870 GND ICV_1 $T=159080 -95435 0 90 $X=158290 $Y=-96095
X1926 361 1120 360 1110 871 GND ICV_1 $T=159080 -89395 0 90 $X=158290 $Y=-90055
X1927 365 1139 364 1127 866 GND ICV_1 $T=163540 -131675 0 90 $X=162750 $Y=-132335
X1928 365 1140 364 1128 867 GND ICV_1 $T=163540 -125635 0 90 $X=162750 $Y=-126295
X1929 365 1141 364 1129 868 GND ICV_1 $T=163540 -119595 0 90 $X=162750 $Y=-120255
X1930 365 1142 364 1130 863 GND ICV_1 $T=163540 -113555 0 90 $X=162750 $Y=-114215
X1931 365 1143 364 1131 864 GND ICV_1 $T=163540 -107515 0 90 $X=162750 $Y=-108175
X1932 365 1144 364 1132 869 GND ICV_1 $T=163540 -101475 0 90 $X=162750 $Y=-102135
X1933 365 1145 364 1133 870 GND ICV_1 $T=163540 -95435 0 90 $X=162750 $Y=-96095
X1934 365 1146 364 1134 871 GND ICV_1 $T=163540 -89395 0 90 $X=162750 $Y=-90055
X1935 369 1163 368 1153 866 GND ICV_1 $T=168000 -131675 0 90 $X=167210 $Y=-132335
X1936 369 1164 368 1154 867 GND ICV_1 $T=168000 -125635 0 90 $X=167210 $Y=-126295
X1937 369 1165 368 1155 868 GND ICV_1 $T=168000 -119595 0 90 $X=167210 $Y=-120255
X1938 369 1166 368 1156 863 GND ICV_1 $T=168000 -113555 0 90 $X=167210 $Y=-114215
X1939 369 1167 368 1157 864 GND ICV_1 $T=168000 -107515 0 90 $X=167210 $Y=-108175
X1940 369 1168 368 1158 869 GND ICV_1 $T=168000 -101475 0 90 $X=167210 $Y=-102135
X1941 369 1169 368 1159 870 GND ICV_1 $T=168000 -95435 0 90 $X=167210 $Y=-96095
X1942 369 1170 368 1160 871 GND ICV_1 $T=168000 -89395 0 90 $X=167210 $Y=-90055
X1943 373 1191 372 1179 866 GND ICV_1 $T=172460 -131675 0 90 $X=171670 $Y=-132335
X1944 373 1192 372 1180 867 GND ICV_1 $T=172460 -125635 0 90 $X=171670 $Y=-126295
X1945 373 1193 372 1181 868 GND ICV_1 $T=172460 -119595 0 90 $X=171670 $Y=-120255
X1946 373 1194 372 1182 863 GND ICV_1 $T=172460 -113555 0 90 $X=171670 $Y=-114215
X1947 373 1195 372 1183 864 GND ICV_1 $T=172460 -107515 0 90 $X=171670 $Y=-108175
X1948 373 1196 372 1184 869 GND ICV_1 $T=172460 -101475 0 90 $X=171670 $Y=-102135
X1949 373 1197 372 1185 870 GND ICV_1 $T=172460 -95435 0 90 $X=171670 $Y=-96095
X1950 373 1198 372 1186 871 GND ICV_1 $T=172460 -89395 0 90 $X=171670 $Y=-90055
X1951 377 1213 376 1203 866 GND ICV_1 $T=176920 -131675 0 90 $X=176130 $Y=-132335
X1952 377 1214 376 1204 867 GND ICV_1 $T=176920 -125635 0 90 $X=176130 $Y=-126295
X1953 377 1215 376 1205 868 GND ICV_1 $T=176920 -119595 0 90 $X=176130 $Y=-120255
X1954 377 1216 376 1206 863 GND ICV_1 $T=176920 -113555 0 90 $X=176130 $Y=-114215
X1955 377 1217 376 1207 864 GND ICV_1 $T=176920 -107515 0 90 $X=176130 $Y=-108175
X1956 377 1218 376 1208 869 GND ICV_1 $T=176920 -101475 0 90 $X=176130 $Y=-102135
X1957 377 1219 376 1209 870 GND ICV_1 $T=176920 -95435 0 90 $X=176130 $Y=-96095
X1958 377 1220 376 1210 871 GND ICV_1 $T=176920 -89395 0 90 $X=176130 $Y=-90055
X1959 381 1241 380 1229 866 GND ICV_1 $T=181380 -131675 0 90 $X=180590 $Y=-132335
X1960 381 1242 380 1230 867 GND ICV_1 $T=181380 -125635 0 90 $X=180590 $Y=-126295
X1961 381 1243 380 1231 868 GND ICV_1 $T=181380 -119595 0 90 $X=180590 $Y=-120255
X1962 381 1244 380 1232 863 GND ICV_1 $T=181380 -113555 0 90 $X=180590 $Y=-114215
X1963 381 1245 380 1233 864 GND ICV_1 $T=181380 -107515 0 90 $X=180590 $Y=-108175
X1964 381 1246 380 1234 869 GND ICV_1 $T=181380 -101475 0 90 $X=180590 $Y=-102135
X1965 381 1247 380 1235 870 GND ICV_1 $T=181380 -95435 0 90 $X=180590 $Y=-96095
X1966 381 1248 380 1236 871 GND ICV_1 $T=181380 -89395 0 90 $X=180590 $Y=-90055
X1967 385 1263 384 1253 866 GND ICV_1 $T=185840 -131675 0 90 $X=185050 $Y=-132335
X1968 385 1264 384 1254 867 GND ICV_1 $T=185840 -125635 0 90 $X=185050 $Y=-126295
X1969 385 1265 384 1255 868 GND ICV_1 $T=185840 -119595 0 90 $X=185050 $Y=-120255
X1970 385 1266 384 1256 863 GND ICV_1 $T=185840 -113555 0 90 $X=185050 $Y=-114215
X1971 385 1267 384 1257 864 GND ICV_1 $T=185840 -107515 0 90 $X=185050 $Y=-108175
X1972 385 1268 384 1258 869 GND ICV_1 $T=185840 -101475 0 90 $X=185050 $Y=-102135
X1973 385 1269 384 1259 870 GND ICV_1 $T=185840 -95435 0 90 $X=185050 $Y=-96095
X1974 385 1270 384 1260 871 GND ICV_1 $T=185840 -89395 0 90 $X=185050 $Y=-90055
X1975 GND 872 324 325 896 897 328 329 922 322 MODE 326 327 330 ICV_3 $T=118450 -154345 0 0 $X=117790 $Y=-155475
X1976 GND 923 332 333 946 947 336 337 972 331 MODE 334 335 338 ICV_3 $T=127370 -154345 0 0 $X=126710 $Y=-155475
X1977 GND 973 340 341 996 999 344 345 1022 339 MODE 342 343 346 ICV_3 $T=136290 -154345 0 0 $X=135630 $Y=-155475
X1978 GND 1023 348 349 1046 1051 352 353 1072 347 MODE 350 351 354 ICV_3 $T=145210 -154345 0 0 $X=144550 $Y=-155475
X1979 GND 1075 356 357 1098 1101 360 361 1122 355 MODE 358 359 362 ICV_3 $T=154130 -154345 0 0 $X=153470 $Y=-155475
X1980 GND 1125 364 365 1150 1151 368 369 1172 363 MODE 366 367 370 ICV_3 $T=163050 -154345 0 0 $X=162390 $Y=-155475
X1981 GND 1175 372 373 1200 1201 376 377 1224 371 MODE 374 375 378 ICV_3 $T=171970 -154345 0 0 $X=171310 $Y=-155475
X1982 GND 1225 380 381 1250 1251 384 385 1272 379 MODE 382 383 386 ICV_3 $T=180890 -154345 0 0 $X=180230 $Y=-155475
X1983 VDD VDD 231 ADD2 p18_CDNS_673890194795 $T=59735 -123355 1 270 $X=58165 $Y=-124445
X1984 VDD VDD 241 ADD1 p18_CDNS_673890194795 $T=59735 -121335 1 270 $X=58165 $Y=-122425
X1985 VDD VDD 234 ADD0 p18_CDNS_673890194795 $T=59735 -119315 1 270 $X=58165 $Y=-120405
X1986 VDD VDD 19 687 p18_CDNS_673890194795 $T=70180 -131555 1 270 $X=68610 $Y=-132645
X1987 VDD VDD 25 688 p18_CDNS_673890194795 $T=70180 -126915 1 270 $X=68610 $Y=-128005
X1988 VDD VDD 24 689 p18_CDNS_673890194795 $T=70180 -122275 1 270 $X=68610 $Y=-123365
X1989 VDD VDD 26 690 p18_CDNS_673890194795 $T=70180 -117635 1 270 $X=68610 $Y=-118725
X1990 VDD VDD 27 691 p18_CDNS_673890194795 $T=70180 -112995 1 270 $X=68610 $Y=-114085
X1991 VDD VDD 21 694 p18_CDNS_673890194795 $T=70180 -99075 1 270 $X=68610 $Y=-100165
X1992 VDD VDD 826 812 p18_CDNS_673890194795 $T=96810 -74465 0 0 $X=95900 $Y=-74895
X1993 VDD VDD 279 275 p18_CDNS_673890194795 $T=101450 -148305 1 0 $X=100540 $Y=-149875
X1994 VDD VDD 292 MODE p18_CDNS_673890194795 $T=105490 -148305 1 0 $X=104580 $Y=-149875
X1995 VDD VDD 859 858 p18_CDNS_673890194795 $T=110810 -150665 0 0 $X=109900 $Y=-151095
X1996 VDD 324 325 328 329 873 ICV_5 $T=118490 -82085 0 0 $X=117580 $Y=-82515
X1997 VDD 332 333 336 337 873 ICV_5 $T=127410 -82085 0 0 $X=126500 $Y=-82515
X1998 VDD 340 341 344 345 873 ICV_5 $T=136330 -82085 0 0 $X=135420 $Y=-82515
X1999 VDD 348 349 352 353 873 ICV_5 $T=145250 -82085 0 0 $X=144340 $Y=-82515
X2000 VDD 356 357 360 361 873 ICV_5 $T=154170 -82085 0 0 $X=153260 $Y=-82515
X2001 VDD 364 365 368 369 873 ICV_5 $T=163090 -82085 0 0 $X=162180 $Y=-82515
X2002 VDD 372 373 376 377 873 ICV_5 $T=172010 -82085 0 0 $X=171100 $Y=-82515
X2003 VDD 380 381 384 385 873 ICV_5 $T=180930 -82085 0 0 $X=180020 $Y=-82515
X2004 VDD 912 39 884 36 GND 921 893 ICV_8 $T=118630 -144565 1 180 $X=117540 $Y=-145695
X2005 VDD 962 43 936 40 GND 971 945 ICV_8 $T=127550 -144565 1 180 $X=126460 $Y=-145695
X2006 VDD 1012 46 986 44 GND 1021 995 ICV_8 $T=136470 -144565 1 180 $X=135380 $Y=-145695
X2007 VDD 1062 51 1036 48 GND 1071 1045 ICV_8 $T=145390 -144565 1 180 $X=144300 $Y=-145695
X2008 VDD 1112 57 1086 55 GND 1121 1097 ICV_8 $T=154310 -144565 1 180 $X=153220 $Y=-145695
X2009 VDD 1162 64 1138 60 GND 1171 1147 ICV_8 $T=163230 -144565 1 180 $X=162140 $Y=-145695
X2010 VDD 1212 69 1190 67 GND 1223 1199 ICV_8 $T=172150 -144565 1 180 $X=171060 $Y=-145695
X2011 VDD 1262 75 1240 72 GND 1271 1249 ICV_8 $T=181070 -144565 1 180 $X=179980 $Y=-145695
X2012 GND VDD 875 885 901 913 925 937 951 963 975 987 1003 1013 1027 1037 1053 1063 1077 1087
+ 1103 1113 1127 1139 1153 1163 1179 1191 1203 1213 1229 1241 1253 1263
+ ICV_15 $T=118450 -130045 0 0 $X=116930 $Y=-130395
X2013 GND VDD 876 886 902 914 926 938 952 964 976 988 1004 1014 1028 1038 1054 1064 1078 1088
+ 1104 1114 1128 1140 1154 1164 1180 1192 1204 1214 1230 1242 1254 1264
+ ICV_15 $T=118450 -124005 0 0 $X=116930 $Y=-124355
X2014 GND VDD 877 887 903 915 927 939 953 965 977 989 1005 1015 1029 1039 1055 1065 1079 1089
+ 1105 1115 1129 1141 1155 1165 1181 1193 1205 1215 1231 1243 1255 1265
+ ICV_15 $T=118450 -117965 0 0 $X=116930 $Y=-118315
X2015 GND VDD 878 888 904 916 928 940 954 966 978 990 1006 1016 1030 1040 1056 1066 1080 1090
+ 1106 1116 1130 1142 1156 1166 1182 1194 1206 1216 1232 1244 1256 1266
+ ICV_15 $T=118450 -111925 0 0 $X=116930 $Y=-112275
X2016 GND VDD 879 889 905 917 929 941 955 967 979 991 1007 1017 1031 1041 1057 1067 1081 1091
+ 1107 1117 1131 1143 1157 1167 1183 1195 1207 1217 1233 1245 1257 1267
+ ICV_15 $T=118450 -105885 0 0 $X=116930 $Y=-106235
X2017 GND VDD 880 890 906 918 930 942 956 968 980 992 1008 1018 1032 1042 1058 1068 1082 1092
+ 1108 1118 1132 1144 1158 1168 1184 1196 1208 1218 1234 1246 1258 1268
+ ICV_15 $T=118450 -99845 0 0 $X=116930 $Y=-100195
X2018 GND VDD 881 891 907 919 931 943 957 969 981 993 1009 1019 1033 1043 1059 1069 1083 1093
+ 1109 1119 1133 1145 1159 1169 1185 1197 1209 1219 1235 1247 1259 1269
+ ICV_15 $T=118450 -93805 0 0 $X=116930 $Y=-94155
X2019 GND VDD 882 892 908 920 932 944 958 970 982 994 1010 1020 1034 1044 1060 1070 1084 1094
+ 1110 1120 1134 1146 1160 1170 1186 1198 1210 1220 1236 1248 1260 1270
+ ICV_15 $T=118450 -87765 0 0 $X=116930 $Y=-88115
X2020 GND 860 859 n18_CDNS_6738901947913 $T=112790 -156365 0 0 $X=112130 $Y=-157495
X2021 GND 323 860 n18_CDNS_6738901947913 $T=114730 -156365 0 0 $X=114070 $Y=-157495
X2022 VDD 860 859 p18_CDNS_6738901947914 $T=112790 -153745 0 0 $X=111880 $Y=-154175
X2023 VDD 323 860 p18_CDNS_6738901947914 $T=114730 -153745 0 0 $X=113820 $Y=-154175
X2024 GND GND 80 78 n18_CDNS_673890194799 $T=-166395 -103525 0 0 $X=-167055 $Y=-104655
X2025 GND GND 84 82 n18_CDNS_673890194799 $T=-155015 -103525 0 0 $X=-155675 $Y=-104655
X2026 GND GND 88 86 n18_CDNS_673890194799 $T=-143635 -103525 0 0 $X=-144295 $Y=-104655
X2027 GND GND 92 90 n18_CDNS_673890194799 $T=-132255 -103525 0 0 $X=-132915 $Y=-104655
X2028 GND GND 96 94 n18_CDNS_673890194799 $T=-120875 -103525 0 0 $X=-121535 $Y=-104655
X2029 GND GND 100 98 n18_CDNS_673890194799 $T=-109495 -103525 0 0 $X=-110155 $Y=-104655
X2030 GND GND 104 102 n18_CDNS_673890194799 $T=-98115 -103525 0 0 $X=-98775 $Y=-104655
X2031 GND GND 108 106 n18_CDNS_673890194799 $T=-86735 -103525 0 0 $X=-87395 $Y=-104655
X2032 GND GND 112 110 n18_CDNS_673890194799 $T=-75355 -103525 0 0 $X=-76015 $Y=-104655
X2033 GND GND 116 114 n18_CDNS_673890194799 $T=-63975 -103525 0 0 $X=-64635 $Y=-104655
X2034 GND GND 120 118 n18_CDNS_673890194799 $T=-52595 -103525 0 0 $X=-53255 $Y=-104655
X2035 GND GND 124 122 n18_CDNS_673890194799 $T=-41215 -103525 0 0 $X=-41875 $Y=-104655
X2036 GND GND 128 126 n18_CDNS_673890194799 $T=-29835 -103525 0 0 $X=-30495 $Y=-104655
X2037 GND GND 132 130 n18_CDNS_673890194799 $T=-18455 -103525 0 0 $X=-19115 $Y=-104655
X2038 GND GND 136 134 n18_CDNS_673890194799 $T=-7075 -103525 0 0 $X=-7735 $Y=-104655
X2039 GND GND 141 138 n18_CDNS_673890194799 $T=4305 -103525 0 0 $X=3645 $Y=-104655
X2040 GND 867 314 MODE n18_CDNS_673890194799 $T=111350 -127365 1 0 $X=110690 $Y=-128155
X2041 GND 868 315 MODE n18_CDNS_673890194799 $T=111350 -125885 0 0 $X=110690 $Y=-127015
X2042 GND 863 316 MODE n18_CDNS_673890194799 $T=111350 -112125 1 0 $X=110690 $Y=-112915
X2043 GND 864 317 MODE n18_CDNS_673890194799 $T=111350 -110645 0 0 $X=110690 $Y=-111775
X2044 GND 869 318 MODE n18_CDNS_673890194799 $T=111350 -96885 1 0 $X=110690 $Y=-97675
X2045 GND 870 319 MODE n18_CDNS_673890194799 $T=111350 -95405 0 0 $X=110690 $Y=-96535
X2046 GND 871 320 MODE n18_CDNS_673890194799 $T=111350 -81645 1 0 $X=110690 $Y=-82435
X2047 GND GND 313 294 n18_CDNS_673890194799 $T=114010 -141125 0 0 $X=113350 $Y=-142255
X2048 GND GND 314 295 n18_CDNS_673890194799 $T=114010 -127365 1 0 $X=113350 $Y=-128155
X2049 GND GND 315 296 n18_CDNS_673890194799 $T=114010 -125885 0 0 $X=113350 $Y=-127015
X2050 GND GND 316 297 n18_CDNS_673890194799 $T=114010 -112125 1 0 $X=113350 $Y=-112915
X2051 GND GND 317 298 n18_CDNS_673890194799 $T=114010 -110645 0 0 $X=113350 $Y=-111775
X2052 GND GND 318 299 n18_CDNS_673890194799 $T=114010 -96885 1 0 $X=113350 $Y=-97675
X2053 GND GND 319 300 n18_CDNS_673890194799 $T=114010 -95405 0 0 $X=113350 $Y=-96535
X2054 GND 861 261 n18_CDNS_6738901947911 $T=112790 -142605 1 0 $X=112130 $Y=-143835
X2055 GND 703 717 698 ICV_16 $T=77370 -80165 0 0 $X=76710 $Y=-81295
X2056 GND 778 790 764 ICV_16 $T=90110 -141125 0 0 $X=89450 $Y=-142255
X2057 GND 275 788 775 ICV_16 $T=90950 -80165 0 0 $X=90290 $Y=-81295
X2058 GND 837 856 827 ICV_16 $T=102250 -156365 0 0 $X=101590 $Y=-157495
X2059 GND 862 873 262 ICV_16 $T=112790 -80165 0 0 $X=112130 $Y=-81295
X2060 VDD 856 837 p18_CDNS_6738901947912 $T=104190 -151985 0 0 $X=103280 $Y=-152415
X2061 VDD 788 812 275 ICV_17 $T=92890 -75785 0 0 $X=91980 $Y=-76215
X2062 VDD 861 865 261 ICV_17 $T=112790 -146985 1 0 $X=111880 $Y=-149875
X2063 VDD 862 873 262 ICV_17 $T=112790 -75785 0 0 $X=111880 $Y=-76215
X2064 VDD MODE 1518 p18_CDNS_673890194794 $T=107470 -147865 1 0 $X=106560 $Y=-149875
X2065 VDD 37 SEL 77 ICV_18 $T=-169055 -98265 0 0 $X=-169965 $Y=-98695
X2066 VDD 38 SEL 81 ICV_18 $T=-157675 -98265 0 0 $X=-158585 $Y=-98695
X2067 VDD 41 SEL 85 ICV_18 $T=-146295 -98265 0 0 $X=-147205 $Y=-98695
X2068 VDD 42 SEL 89 ICV_18 $T=-134915 -98265 0 0 $X=-135825 $Y=-98695
X2069 VDD 45 SEL 93 ICV_18 $T=-123535 -98265 0 0 $X=-124445 $Y=-98695
X2070 VDD 47 SEL 97 ICV_18 $T=-112155 -98265 0 0 $X=-113065 $Y=-98695
X2071 VDD 49 SEL 101 ICV_18 $T=-100775 -98265 0 0 $X=-101685 $Y=-98695
X2072 VDD 52 SEL 105 ICV_18 $T=-89395 -98265 0 0 $X=-90305 $Y=-98695
X2073 VDD 56 SEL 109 ICV_18 $T=-78015 -98265 0 0 $X=-78925 $Y=-98695
X2074 VDD 58 SEL 113 ICV_18 $T=-66635 -98265 0 0 $X=-67545 $Y=-98695
X2075 VDD 62 SEL 117 ICV_18 $T=-55255 -98265 0 0 $X=-56165 $Y=-98695
X2076 VDD 66 SEL 121 ICV_18 $T=-43875 -98265 0 0 $X=-44785 $Y=-98695
X2077 VDD 68 SEL 125 ICV_18 $T=-32495 -98265 0 0 $X=-33405 $Y=-98695
X2078 VDD 71 SEL 129 ICV_18 $T=-21115 -98265 0 0 $X=-22025 $Y=-98695
X2079 VDD 74 SEL 133 ICV_18 $T=-9735 -98265 0 0 $X=-10645 $Y=-98695
X2080 VDD 76 SEL 137 ICV_18 $T=1645 -98265 0 0 $X=735 $Y=-98695
X2081 VDD 262 MODE 280 ICV_18 $T=107470 -74905 0 0 $X=106560 $Y=-75335
X2082 VDD 866 MODE 284 ICV_18 $T=111350 -135865 0 0 $X=110440 $Y=-136295
X2083 VDD 867 MODE 285 ICV_18 $T=111350 -132625 1 0 $X=110440 $Y=-134635
X2084 VDD 868 MODE 286 ICV_18 $T=111350 -120625 0 0 $X=110440 $Y=-121055
X2085 VDD 863 MODE 287 ICV_18 $T=111350 -117385 1 0 $X=110440 $Y=-119395
X2086 VDD 864 MODE 288 ICV_18 $T=111350 -105385 0 0 $X=110440 $Y=-105815
X2087 VDD 869 MODE 289 ICV_18 $T=111350 -102145 1 0 $X=110440 $Y=-104155
X2088 VDD 870 MODE 290 ICV_18 $T=111350 -90145 0 0 $X=110440 $Y=-90575
X2089 VDD 871 MODE 291 ICV_18 $T=111350 -86905 1 0 $X=110440 $Y=-88915
X2090 GND 798 790 n18_CDNS_673890194798 $T=94030 -141025 0 0 $X=93330 $Y=-142255
X2091 GND 805 797 n18_CDNS_673890194798 $T=94030 -81745 1 0 $X=93330 $Y=-82315
X2092 GND 826 812 n18_CDNS_673890194798 $T=96810 -80065 0 0 $X=96110 $Y=-81295
X2093 GND 828 817 n18_CDNS_673890194798 $T=98670 -141025 0 0 $X=97970 $Y=-142255
X2094 GND 835 824 n18_CDNS_673890194798 $T=98670 -81745 1 0 $X=97970 $Y=-82315
X2095 GND 293 MODE n18_CDNS_673890194798 $T=105490 -80065 0 0 $X=104790 $Y=-81295
X2096 GND 857 856 n18_CDNS_673890194798 $T=106170 -156265 0 0 $X=105470 $Y=-157495
X2097 GND 859 858 n18_CDNS_673890194798 $T=110810 -156265 0 0 $X=110110 $Y=-157495
X2098 GND 866 313 305 MODE ICV_19 $T=109370 -141025 0 0 $X=108670 $Y=-142255
X2099 GND 817 264 1394 n18_CDNS_673890194797 $T=96440 -141125 0 0 $X=96120 $Y=-142255
X2100 GND 818 265 1395 n18_CDNS_673890194797 $T=96440 -127365 1 0 $X=96120 $Y=-128155
X2101 GND 819 266 1396 n18_CDNS_673890194797 $T=96440 -125885 0 0 $X=96120 $Y=-127015
X2102 GND 820 267 1397 n18_CDNS_673890194797 $T=96440 -112125 1 0 $X=96120 $Y=-112915
X2103 GND 821 268 1398 n18_CDNS_673890194797 $T=96440 -110645 0 0 $X=96120 $Y=-111775
X2104 GND 822 269 1399 n18_CDNS_673890194797 $T=96440 -96885 1 0 $X=96120 $Y=-97675
X2105 GND 823 270 1400 n18_CDNS_673890194797 $T=96440 -95405 0 0 $X=96120 $Y=-96535
X2106 GND 839 829 1401 n18_CDNS_673890194797 $T=101080 -127365 1 0 $X=100760 $Y=-128155
X2107 GND 840 830 1402 n18_CDNS_673890194797 $T=101080 -125885 0 0 $X=100760 $Y=-127015
X2108 GND 841 831 1403 n18_CDNS_673890194797 $T=101080 -112125 1 0 $X=100760 $Y=-112915
X2109 GND 842 832 1404 n18_CDNS_673890194797 $T=101080 -110645 0 0 $X=100760 $Y=-111775
X2110 GND 843 833 1405 n18_CDNS_673890194797 $T=101080 -96885 1 0 $X=100760 $Y=-97675
X2111 GND 844 834 1406 n18_CDNS_673890194797 $T=101080 -95405 0 0 $X=100760 $Y=-96535
X2112 GND 858 857 1407 n18_CDNS_673890194797 $T=108580 -156365 0 0 $X=108260 $Y=-157495
X2113 GND 798 1394 n18_CDNS_673890194796 $T=96010 -141125 0 0 $X=95350 $Y=-142255
X2114 GND 799 1395 n18_CDNS_673890194796 $T=96010 -127365 1 0 $X=95350 $Y=-128155
X2115 GND 800 1396 n18_CDNS_673890194796 $T=96010 -125885 0 0 $X=95350 $Y=-127015
X2116 GND 801 1397 n18_CDNS_673890194796 $T=96010 -112125 1 0 $X=95350 $Y=-112915
X2117 GND 802 1398 n18_CDNS_673890194796 $T=96010 -110645 0 0 $X=95350 $Y=-111775
X2118 GND 803 1399 n18_CDNS_673890194796 $T=96010 -96885 1 0 $X=95350 $Y=-97675
X2119 GND 804 1400 n18_CDNS_673890194796 $T=96010 -95405 0 0 $X=95350 $Y=-96535
X2120 GND 805 1356 n18_CDNS_673890194796 $T=96010 -81645 1 0 $X=95350 $Y=-82435
X2121 GND 19 1360 n18_CDNS_673890194796 $T=100650 -141125 0 0 $X=99990 $Y=-142255
X2122 GND 25 1401 n18_CDNS_673890194796 $T=100650 -127365 1 0 $X=99990 $Y=-128155
X2123 GND 24 1402 n18_CDNS_673890194796 $T=100650 -125885 0 0 $X=99990 $Y=-127015
X2124 GND 26 1403 n18_CDNS_673890194796 $T=100650 -112125 1 0 $X=99990 $Y=-112915
X2125 GND 27 1404 n18_CDNS_673890194796 $T=100650 -110645 0 0 $X=99990 $Y=-111775
X2126 GND 23 1405 n18_CDNS_673890194796 $T=100650 -96885 1 0 $X=99990 $Y=-97675
X2127 GND 22 1406 n18_CDNS_673890194796 $T=100650 -95405 0 0 $X=99990 $Y=-96535
X2128 GND 21 1361 n18_CDNS_673890194796 $T=100650 -81645 1 0 $X=99990 $Y=-82435
X2129 GND 304 1407 n18_CDNS_673890194796 $T=108150 -156365 0 0 $X=107490 $Y=-157495
X2130 VDD 687 CLK p18_CDNS_673890194790 $T=70620 -128895 1 270 $X=68610 $Y=-129985
X2131 VDD 688 CLK p18_CDNS_673890194790 $T=70620 -124255 1 270 $X=68610 $Y=-125345
X2132 VDD 689 CLK p18_CDNS_673890194790 $T=70620 -119615 1 270 $X=68610 $Y=-120705
X2133 VDD 690 CLK p18_CDNS_673890194790 $T=70620 -114975 1 270 $X=68610 $Y=-116065
X2134 VDD 691 CLK p18_CDNS_673890194790 $T=70620 -110335 1 270 $X=68610 $Y=-111425
X2135 VDD 692 CLK p18_CDNS_673890194790 $T=70620 -105695 1 270 $X=68610 $Y=-106785
X2136 VDD 836 CLK p18_CDNS_673890194790 $T=98790 -74905 0 0 $X=97880 $Y=-75335
X2137 VDD 858 304 p18_CDNS_673890194790 $T=108150 -151105 0 0 $X=107240 $Y=-151535
X2138 GND 708 264 262 708 ICV_20 $T=78350 -141025 0 0 $X=77650 $Y=-142255
X2139 GND 280 282 836 VDD ICV_20 $T=101450 -80065 0 0 $X=100750 $Y=-81295
X2140 GND 301 312 21 MODE ICV_20 $T=107350 -81745 1 0 $X=106650 $Y=-82315
X2141 GND 800 799 792 791 ICV_21 $T=94030 -127465 1 0 $X=93330 $Y=-128035
X2142 GND 802 801 794 793 ICV_21 $T=94030 -112225 1 0 $X=93330 $Y=-112795
X2143 GND 804 803 796 795 ICV_21 $T=94030 -96985 1 0 $X=93330 $Y=-97555
X2144 GND 830 829 819 818 ICV_21 $T=98670 -127465 1 0 $X=97970 $Y=-128035
X2145 GND 832 831 821 820 ICV_21 $T=98670 -112225 1 0 $X=97970 $Y=-112795
X2146 GND 834 833 823 822 ICV_21 $T=98670 -96985 1 0 $X=97970 $Y=-97555
X2147 GND 710 709 266 265 262 262 710 709 ICV_22 $T=78350 -127465 1 0 $X=77650 $Y=-128035
X2148 GND 712 711 268 267 262 262 712 711 ICV_22 $T=78350 -112225 1 0 $X=77650 $Y=-112795
X2149 GND 714 713 270 269 262 262 714 713 ICV_22 $T=78350 -96985 1 0 $X=77650 $Y=-97555
X2150 GND 850 849 286 285 840 839 850 849 ICV_22 $T=103310 -127465 1 0 $X=102610 $Y=-128035
X2151 GND 852 851 288 287 842 841 852 851 ICV_22 $T=103310 -112225 1 0 $X=102610 $Y=-112795
X2152 GND 854 853 290 289 844 843 854 853 ICV_22 $T=103310 -96985 1 0 $X=102610 $Y=-97555
X2153 GND 296 295 307 306 24 25 MODE MODE ICV_22 $T=107350 -127465 1 0 $X=106650 $Y=-128035
X2154 GND 298 297 309 308 27 26 MODE MODE ICV_22 $T=107350 -112225 1 0 $X=106650 $Y=-112795
X2155 GND 300 299 311 310 22 23 MODE MODE ICV_22 $T=107350 -96985 1 0 $X=106650 $Y=-97555
X2156 VDD 798 799 790 791 ICV_23 $T=94030 -135425 0 0 $X=93120 $Y=-135855
X2157 VDD 800 801 792 793 ICV_23 $T=94030 -120185 0 0 $X=93120 $Y=-120615
X2158 VDD 802 803 794 795 ICV_23 $T=94030 -104945 0 0 $X=93120 $Y=-105375
X2159 VDD 804 805 796 797 ICV_23 $T=94030 -89705 0 0 $X=93120 $Y=-90135
X2160 VDD 828 829 817 818 ICV_23 $T=98670 -135425 0 0 $X=97760 $Y=-135855
X2161 VDD 830 831 819 820 ICV_23 $T=98670 -120185 0 0 $X=97760 $Y=-120615
X2162 VDD 832 833 821 822 ICV_23 $T=98670 -104945 0 0 $X=97760 $Y=-105375
X2163 VDD 834 835 823 824 ICV_23 $T=98670 -89705 0 0 $X=97760 $Y=-90135
X2164 VDD 708 709 264 265 262 262 708 709 ICV_24 $T=78350 -135425 0 0 $X=77440 $Y=-135855
X2165 VDD 710 711 266 267 262 262 710 711 ICV_24 $T=78350 -120185 0 0 $X=77440 $Y=-120615
X2166 VDD 712 713 268 269 262 262 712 713 ICV_24 $T=78350 -104945 0 0 $X=77440 $Y=-105375
X2167 VDD 714 715 270 271 262 262 714 715 ICV_24 $T=78350 -89705 0 0 $X=77440 $Y=-90135
X2168 VDD 848 849 284 285 838 839 848 849 ICV_24 $T=103310 -135425 0 0 $X=102400 $Y=-135855
X2169 VDD 850 851 286 287 840 841 850 851 ICV_24 $T=103310 -120185 0 0 $X=102400 $Y=-120615
X2170 VDD 852 853 288 289 842 843 852 853 ICV_24 $T=103310 -104945 0 0 $X=102400 $Y=-105375
X2171 VDD 854 855 290 291 844 845 854 855 ICV_24 $T=103310 -89705 0 0 $X=102400 $Y=-90135
X2172 VDD 294 295 305 306 19 25 MODE MODE ICV_24 $T=107350 -135425 0 0 $X=106440 $Y=-135855
X2173 VDD 296 297 307 308 24 26 MODE MODE ICV_24 $T=107350 -120185 0 0 $X=106440 $Y=-120615
X2174 VDD 298 299 309 310 27 23 MODE MODE ICV_24 $T=107350 -104945 0 0 $X=106440 $Y=-105375
X2175 VDD 300 301 311 312 22 21 MODE MODE ICV_24 $T=107350 -89705 0 0 $X=106440 $Y=-90135
X2176 GND 79 37 80 77 78 SEL IN0 Q0 ICV_25 $T=-175075 -103425 0 0 $X=-175775 $Y=-104655
X2177 GND 83 38 84 81 82 SEL IN1 Q1 ICV_25 $T=-163695 -103425 0 0 $X=-164395 $Y=-104655
X2178 GND 87 41 88 85 86 SEL IN2 Q2 ICV_25 $T=-152315 -103425 0 0 $X=-153015 $Y=-104655
X2179 GND 91 42 92 89 90 SEL IN3 Q3 ICV_25 $T=-140935 -103425 0 0 $X=-141635 $Y=-104655
X2180 GND 95 45 96 93 94 SEL IN4 Q4 ICV_25 $T=-129555 -103425 0 0 $X=-130255 $Y=-104655
X2181 GND 99 47 100 97 98 SEL IN5 Q5 ICV_25 $T=-118175 -103425 0 0 $X=-118875 $Y=-104655
X2182 GND 103 49 104 101 102 SEL IN6 Q6 ICV_25 $T=-106795 -103425 0 0 $X=-107495 $Y=-104655
X2183 GND 107 52 108 105 106 SEL IN7 Q7 ICV_25 $T=-95415 -103425 0 0 $X=-96115 $Y=-104655
X2184 GND 111 56 112 109 110 SEL IN8 Q8 ICV_25 $T=-84035 -103425 0 0 $X=-84735 $Y=-104655
X2185 GND 115 58 116 113 114 SEL IN9 GND ICV_25 $T=-72655 -103425 0 0 $X=-73355 $Y=-104655
X2186 GND 119 62 120 117 118 SEL IN10 GND ICV_25 $T=-61275 -103425 0 0 $X=-61975 $Y=-104655
X2187 GND 123 66 124 121 122 SEL IN11 GND ICV_25 $T=-49895 -103425 0 0 $X=-50595 $Y=-104655
X2188 GND 127 68 128 125 126 SEL IN12 GND ICV_25 $T=-38515 -103425 0 0 $X=-39215 $Y=-104655
X2189 GND 131 71 132 129 130 SEL IN13 GND ICV_25 $T=-27135 -103425 0 0 $X=-27835 $Y=-104655
X2190 GND 135 74 136 133 134 SEL IN14 GND ICV_25 $T=-15755 -103425 0 0 $X=-16455 $Y=-104655
X2191 GND 140 76 141 137 138 SEL IN15 GND ICV_25 $T=-4375 -103425 0 0 $X=-5075 $Y=-104655
X2192 GND 292 261 302 279 281 MODE 275 GND ICV_25 $T=101450 -142705 1 0 $X=100750 $Y=-143395
X2193 VDD 77 78 79 IN0 Q0 SEL ICV_26 $T=-175075 -97825 0 0 $X=-175985 $Y=-98255
X2194 VDD 81 82 83 IN1 Q1 SEL ICV_26 $T=-163695 -97825 0 0 $X=-164605 $Y=-98255
X2195 VDD 85 86 87 IN2 Q2 SEL ICV_26 $T=-152315 -97825 0 0 $X=-153225 $Y=-98255
X2196 VDD 89 90 91 IN3 Q3 SEL ICV_26 $T=-140935 -97825 0 0 $X=-141845 $Y=-98255
X2197 VDD 93 94 95 IN4 Q4 SEL ICV_26 $T=-129555 -97825 0 0 $X=-130465 $Y=-98255
X2198 VDD 97 98 99 IN5 Q5 SEL ICV_26 $T=-118175 -97825 0 0 $X=-119085 $Y=-98255
X2199 VDD 101 102 103 IN6 Q6 SEL ICV_26 $T=-106795 -97825 0 0 $X=-107705 $Y=-98255
X2200 VDD 105 106 107 IN7 Q7 SEL ICV_26 $T=-95415 -97825 0 0 $X=-96325 $Y=-98255
X2201 VDD 109 110 111 IN8 Q8 SEL ICV_26 $T=-84035 -97825 0 0 $X=-84945 $Y=-98255
X2202 VDD 113 114 115 IN9 GND SEL ICV_26 $T=-72655 -97825 0 0 $X=-73565 $Y=-98255
X2203 VDD 117 118 119 IN10 GND SEL ICV_26 $T=-61275 -97825 0 0 $X=-62185 $Y=-98255
X2204 VDD 121 122 123 IN11 GND SEL ICV_26 $T=-49895 -97825 0 0 $X=-50805 $Y=-98255
X2205 VDD 125 126 127 IN12 GND SEL ICV_26 $T=-38515 -97825 0 0 $X=-39425 $Y=-98255
X2206 VDD 129 130 131 IN13 GND SEL ICV_26 $T=-27135 -97825 0 0 $X=-28045 $Y=-98255
X2207 VDD 133 134 135 IN14 GND SEL ICV_26 $T=-15755 -97825 0 0 $X=-16665 $Y=-98255
X2208 VDD 137 138 140 IN15 GND SEL ICV_26 $T=-4375 -97825 0 0 $X=-5285 $Y=-98255
X2209 VDD 280 282 293 836 VDD MODE ICV_26 $T=101450 -74465 0 0 $X=100540 $Y=-74895
X2210 VDD 817 818 798 799 ICV_27 $T=96010 -135865 0 0 $X=95100 $Y=-136295
X2211 VDD 819 820 800 801 ICV_27 $T=96010 -120625 0 0 $X=95100 $Y=-121055
X2212 VDD 821 822 802 803 ICV_27 $T=96010 -105385 0 0 $X=95100 $Y=-105815
X2213 VDD 823 824 804 805 ICV_27 $T=96010 -90145 0 0 $X=95100 $Y=-90575
X2214 VDD 838 839 19 25 ICV_27 $T=100650 -135865 0 0 $X=99740 $Y=-136295
X2215 VDD 840 841 24 26 ICV_27 $T=100650 -120625 0 0 $X=99740 $Y=-121055
X2216 VDD 842 843 27 23 ICV_27 $T=100650 -105385 0 0 $X=99740 $Y=-105815
X2217 VDD 844 845 22 21 ICV_27 $T=100650 -90145 0 0 $X=99740 $Y=-90575
X2218 GND 724 723 738 737 266 265 ICV_29 $T=82350 -127365 1 0 $X=81690 $Y=-128595
X2219 GND 726 725 740 739 268 267 ICV_29 $T=82350 -112125 1 0 $X=81690 $Y=-113355
X2220 GND 728 727 742 741 270 269 ICV_29 $T=82350 -96885 1 0 $X=81690 $Y=-98115
X2221 GND 752 751 766 765 738 737 ICV_29 $T=86230 -127365 1 0 $X=85570 $Y=-128595
X2222 GND 754 753 768 767 740 739 ICV_29 $T=86230 -112125 1 0 $X=85570 $Y=-113355
X2223 GND 756 755 770 769 742 741 ICV_29 $T=86230 -96885 1 0 $X=85570 $Y=-98115
X2224 GND 780 779 792 791 766 765 ICV_29 $T=90110 -127365 1 0 $X=89450 $Y=-128595
X2225 GND 782 781 794 793 768 767 ICV_29 $T=90110 -112125 1 0 $X=89450 $Y=-113355
X2226 GND 784 783 796 795 770 769 ICV_29 $T=90110 -96885 1 0 $X=89450 $Y=-98115
X2227 VDD 778 790 779 791 764 765 ICV_30 $T=90110 -136745 0 0 $X=89200 $Y=-137175
X2228 VDD 780 792 781 793 766 767 ICV_30 $T=90110 -121505 0 0 $X=89200 $Y=-121935
X2229 VDD 782 794 783 795 768 769 ICV_30 $T=90110 -106265 0 0 $X=89200 $Y=-106695
X2230 VDD 784 796 785 797 770 771 ICV_30 $T=90110 -91025 0 0 $X=89200 $Y=-91455
X2231 GND 722 736 750 764 264 ICV_31 $T=82350 -141125 0 0 $X=81690 $Y=-142255
X2232 GND 733 747 759 775 719 ICV_31 $T=83190 -80165 0 0 $X=82530 $Y=-81295
X2233 GND 448 453 470 485 500 511 516 523 261 ICV_32 $T=24650 -156365 0 0 $X=23990 $Y=-157495
X2234 GND 536 549 556 569 576 585 598 607 523 ICV_32 $T=40170 -156365 0 0 $X=39510 $Y=-157495
X2235 GND 614 617 630 643 651 657 663 669 607 ICV_32 $T=55690 -156365 0 0 $X=55030 $Y=-157495
X2236 GND 644 656 660 668 672 682 686 698 CLK ICV_32 $T=61850 -80165 0 0 $X=61190 $Y=-81295
X2237 GND 681 685 697 304 716 718 730 744 669 ICV_32 $T=71210 -156365 0 0 $X=70550 $Y=-157495
X2238 GND 758 773 786 787 809 814 825 827 744 ICV_32 $T=86730 -156365 0 0 $X=86070 $Y=-157495
X2239 VDD 448 453 470 485 500 511 516 523 261 ICV_34 $T=24650 -151985 0 0 $X=23740 $Y=-152415
X2240 VDD 536 549 556 569 576 585 598 607 523 ICV_34 $T=40170 -151985 0 0 $X=39260 $Y=-152415
X2241 VDD 614 617 630 643 651 657 663 669 607 ICV_34 $T=55690 -151985 0 0 $X=54780 $Y=-152415
X2242 VDD 644 656 660 668 672 682 686 698 CLK ICV_34 $T=61850 -75785 0 0 $X=60940 $Y=-76215
X2243 VDD 681 685 697 304 716 718 730 744 669 ICV_34 $T=71210 -151985 0 0 $X=70300 $Y=-152415
X2244 VDD 703 717 719 733 747 759 775 275 698 ICV_34 $T=77370 -75785 0 0 $X=76460 $Y=-76215
X2245 VDD 758 773 786 787 809 814 825 827 744 ICV_34 $T=86730 -151985 0 0 $X=85820 $Y=-152415
X2246 VDD 722 723 736 737 750 751 764 765 264 265 ICV_35 $T=82350 -136745 0 0 $X=81440 $Y=-137175
X2247 VDD 724 725 738 739 752 753 766 767 266 267 ICV_35 $T=82350 -121505 0 0 $X=81440 $Y=-121935
X2248 VDD 726 727 740 741 754 755 768 769 268 269 ICV_35 $T=82350 -106265 0 0 $X=81440 $Y=-106695
X2249 VDD 728 729 742 743 756 757 770 771 270 271 ICV_35 $T=82350 -91025 0 0 $X=81440 $Y=-91455
X2250 GND 19 687 247 CLK ICV_36 $T=75780 -131555 1 270 $X=75090 $Y=-132435
X2251 GND 25 688 253 CLK ICV_36 $T=75780 -126915 1 270 $X=75090 $Y=-127795
X2252 GND 24 689 254 CLK ICV_36 $T=75780 -122275 1 270 $X=75090 $Y=-123155
X2253 GND 26 690 255 CLK ICV_36 $T=75780 -117635 1 270 $X=75090 $Y=-118515
X2254 GND 27 691 256 CLK ICV_36 $T=75780 -112995 1 270 $X=75090 $Y=-113875
X2255 GND 23 692 257 CLK ICV_36 $T=75780 -108355 1 270 $X=75090 $Y=-109235
X2256 GND 22 693 248 CLK ICV_36 $T=75780 -103715 1 270 $X=75090 $Y=-104595
X2257 GND 21 694 249 CLK ICV_36 $T=75780 -99075 1 270 $X=75090 $Y=-99955
X2258 VDD 234 1561 p18_CDNS_673890194791 $T=66940 -107275 0 270 $X=66510 $Y=-108010
X2259 VDD ADD0 1562 p18_CDNS_673890194791 $T=66940 -103655 0 270 $X=66510 $Y=-104390
X2260 VDD 234 1494 p18_CDNS_673890194791 $T=66940 -100035 0 270 $X=66510 $Y=-100770
X2261 VDD ADD0 1563 p18_CDNS_673890194791 $T=66940 -96415 0 270 $X=66510 $Y=-97150
X2262 VDD 241 1487 1486 p18_CDNS_673890194792 $T=66940 -122185 0 270 $X=66510 $Y=-122920
X2263 VDD ADD1 1492 1564 p18_CDNS_673890194792 $T=66940 -111325 0 270 $X=66510 $Y=-112060
X2264 VDD 241 1561 1565 p18_CDNS_673890194792 $T=66940 -107705 0 270 $X=66510 $Y=-108440
X2265 VDD 241 1562 1566 p18_CDNS_673890194792 $T=66940 -104085 0 270 $X=66510 $Y=-104820
X2266 VDD ADD1 1563 1567 p18_CDNS_673890194792 $T=66940 -96845 0 270 $X=66510 $Y=-97580
X2267 VDD 255 231 1564 p18_CDNS_673890194793 $T=66940 -111755 0 270 $X=66510 $Y=-112845
X2268 VDD 256 ADD2 1565 p18_CDNS_673890194793 $T=66940 -108135 0 270 $X=66510 $Y=-109225
X2269 VDD 257 ADD2 1566 p18_CDNS_673890194793 $T=66940 -104515 0 270 $X=66510 $Y=-105605
X2270 VDD 248 ADD2 1493 p18_CDNS_673890194793 $T=66940 -100895 0 270 $X=66510 $Y=-101985
X2271 VDD 249 ADD2 1567 p18_CDNS_673890194793 $T=66940 -97275 0 270 $X=66510 $Y=-98365
X2272 GND GND 231 ADD2 n18_CDNS_6738901947927 $T=63270 -123355 1 270 $X=62700 $Y=-124235
X2273 GND GND 241 ADD1 n18_CDNS_6738901947927 $T=63270 -121335 1 270 $X=62700 $Y=-122215
X2274 GND 247 GND 231 n18_CDNS_6738901947927 $T=64770 -123355 0 270 $X=63630 $Y=-124235
X2275 GND 253 GND ADD0 n18_CDNS_6738901947927 $T=64770 -118135 0 270 $X=63630 $Y=-119015
X2276 GND 254 GND 231 n18_CDNS_6738901947927 $T=64770 -116115 0 270 $X=63630 $Y=-116995
X2277 GND 254 GND 234 n18_CDNS_6738901947927 $T=64770 -114515 0 270 $X=63630 $Y=-115395
X2278 GND 255 GND 231 n18_CDNS_6738901947927 $T=64770 -112495 0 270 $X=63630 $Y=-113375
X2279 GND 255 GND ADD0 n18_CDNS_6738901947927 $T=64770 -110895 0 270 $X=63630 $Y=-111775
X2280 GND 256 GND ADD2 n18_CDNS_6738901947927 $T=64770 -108875 0 270 $X=63630 $Y=-109755
X2281 GND 256 GND 234 n18_CDNS_6738901947927 $T=64770 -107275 0 270 $X=63630 $Y=-108155
X2282 GND 257 GND ADD2 n18_CDNS_6738901947927 $T=64770 -105255 0 270 $X=63630 $Y=-106135
X2283 GND 257 GND ADD0 n18_CDNS_6738901947927 $T=64770 -103655 0 270 $X=63630 $Y=-104535
X2284 GND 248 GND ADD2 n18_CDNS_6738901947927 $T=64770 -101635 0 270 $X=63630 $Y=-102515
X2285 GND 248 GND 234 n18_CDNS_6738901947927 $T=64770 -100035 0 270 $X=63630 $Y=-100915
X2286 GND 249 GND ADD2 n18_CDNS_6738901947927 $T=64770 -98015 0 270 $X=63630 $Y=-98895
X2287 GND 249 GND ADD0 n18_CDNS_6738901947927 $T=64770 -96415 0 270 $X=63630 $Y=-97295
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT MA C CIN A B GND VDD S
** N=19 EP=7 IP=0 FDC=28
M0 GND 5 C GND NM L=1.8e-07 W=4.4e-07 $X=28980 $Y=-20560 $D=0
M1 GND A 2 GND NM L=1.8e-07 W=4.4e-07 $X=30920 $Y=-20560 $D=0
M2 14 A GND GND NM L=1.8e-07 W=4.4e-07 $X=31640 $Y=-20560 $D=0
M3 5 B 14 GND NM L=1.8e-07 W=4.4e-07 $X=32070 $Y=-20560 $D=0
M4 2 CIN 5 GND NM L=1.8e-07 W=4.4e-07 $X=32790 $Y=-20560 $D=0
M5 GND B 2 GND NM L=1.8e-07 W=4.4e-07 $X=33510 $Y=-20560 $D=0
M6 15 B GND GND NM L=1.8e-07 W=4.4e-07 $X=34230 $Y=-20560 $D=0
M7 16 A 15 GND NM L=1.8e-07 W=4.4e-07 $X=34660 $Y=-20560 $D=0
M8 10 CIN 16 GND NM L=1.8e-07 W=4.4e-07 $X=35090 $Y=-20560 $D=0
M9 7 5 10 GND NM L=1.8e-07 W=4.4e-07 $X=35810 $Y=-20560 $D=0
M10 GND CIN 7 GND NM L=1.8e-07 W=4.4e-07 $X=36530 $Y=-20560 $D=0
M11 7 A GND GND NM L=1.8e-07 W=4.4e-07 $X=37250 $Y=-20560 $D=0
M12 GND B 7 GND NM L=1.8e-07 W=4.4e-07 $X=37970 $Y=-20560 $D=0
M13 S 10 GND GND NM L=1.8e-07 W=4.4e-07 $X=38690 $Y=-20560 $D=0
M14 VDD 5 C VDD PM L=1.8e-07 W=8.8e-07 $X=28980 $Y=-17555 $D=4
M15 VDD A 3 VDD PM L=1.8e-07 W=8.8e-07 $X=30920 $Y=-17555 $D=4
M16 17 A VDD VDD PM L=1.8e-07 W=8.8e-07 $X=31640 $Y=-17555 $D=4
M17 5 B 17 VDD PM L=1.8e-07 W=8.8e-07 $X=32070 $Y=-17555 $D=4
M18 3 CIN 5 VDD PM L=1.8e-07 W=8.8e-07 $X=32790 $Y=-17555 $D=4
M19 VDD B 3 VDD PM L=1.8e-07 W=8.8e-07 $X=33510 $Y=-17555 $D=4
M20 18 B VDD VDD PM L=1.8e-07 W=8.8e-07 $X=34230 $Y=-17555 $D=4
M21 19 A 18 VDD PM L=1.8e-07 W=8.8e-07 $X=34660 $Y=-17555 $D=4
M22 10 CIN 19 VDD PM L=1.8e-07 W=8.8e-07 $X=35090 $Y=-17555 $D=4
M23 8 5 10 VDD PM L=1.8e-07 W=8.8e-07 $X=35810 $Y=-17555 $D=4
M24 VDD CIN 8 VDD PM L=1.8e-07 W=8.8e-07 $X=36530 $Y=-17555 $D=4
M25 8 A VDD VDD PM L=1.8e-07 W=8.8e-07 $X=37250 $Y=-17555 $D=4
M26 VDD B 8 VDD PM L=1.8e-07 W=8.8e-07 $X=37970 $Y=-17555 $D=4
M27 S 10 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=38690 $Y=-17555 $D=4
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_672673910980 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_672673910984 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_672673910983 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672673910981 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 4 3 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672673910982 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT CSA_C COUT B A S INVCI CI VDD GND
** N=22 EP=8 IP=63 FDC=36
M0 8 CI COUT GND NM L=1.8e-07 W=4.4e-07 $X=-1755 $Y=-16485 $D=0
M1 GND 9 8 GND NM L=1.8e-07 W=4.4e-07 $X=-1035 $Y=-16485 $D=0
M2 GND 10 7 GND NM L=1.8e-07 W=4.4e-07 $X=-835 $Y=-12785 $D=0
M3 9 A GND GND NM L=1.8e-07 W=2.2e-07 $X=-275 $Y=-16385 $D=0
M4 19 B GND GND NM L=1.8e-07 W=4.4e-07 $X=-115 $Y=-12785 $D=0
M5 10 A 19 GND NM L=1.8e-07 W=4.4e-07 $X=315 $Y=-12785 $D=0
M6 GND B 9 GND NM L=1.8e-07 W=2.2e-07 $X=525 $Y=-16385 $D=0
M7 13 10 11 GND NM L=1.8e-07 W=4.4e-07 $X=2255 $Y=-12785 $D=0
M8 20 A 14 GND NM L=1.8e-07 W=4.4e-07 $X=2505 $Y=-16485 $D=0
M9 GND B 20 GND NM L=1.8e-07 W=4.4e-07 $X=2935 $Y=-16485 $D=0
M10 GND B 13 GND NM L=1.8e-07 W=4.4e-07 $X=2975 $Y=-12785 $D=0
M11 14 9 GND GND NM L=1.8e-07 W=2.2e-07 $X=3695 $Y=-16385 $D=0
M12 13 A GND GND NM L=1.8e-07 W=4.4e-07 $X=3695 $Y=-12785 $D=0
M13 17 14 GND GND NM L=1.8e-07 W=4.4e-07 $X=5675 $Y=-16485 $D=0
M14 18 11 GND GND NM L=1.8e-07 W=4.4e-07 $X=5675 $Y=-12785 $D=0
M15 S CI 17 GND NM L=1.8e-07 W=4.4e-07 $X=6435 $Y=-16485 $D=0
M16 7 CI COUT VDD PM L=1.8e-07 W=4.4e-07 $X=-1635 $Y=-9340 $D=4
M17 VDD 9 8 VDD PM L=1.8e-07 W=8.8e-07 $X=-835 $Y=-19930 $D=4
M18 10 B VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-115 $Y=-9340 $D=4
M19 11 10 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=2545 $Y=-9340 $D=4
M20 12 B VDD VDD PM L=1.8e-07 W=8.8e-07 $X=2975 $Y=-19930 $D=4
M21 S INVCI 17 VDD PM L=1.8e-07 W=4.4e-07 $X=6395 $Y=-19930 $D=4
M22 S CI 18 VDD PM L=1.8e-07 W=4.4e-07 $X=6435 $Y=-9340 $D=4
X23 VDD 8 COUT INVCI p18_CDNS_672673910980 $T=-1415 -19490 0 180 $X=-2505 $Y=-21280
X24 VDD 10 VDD A p18_CDNS_672673910980 $T=605 -9340 0 0 $X=-305 $Y=-9770
X25 GND 7 COUT INVCI n18_CDNS_672673910984 $T=-1455 -12785 1 180 $X=-2295 $Y=-14805
X26 GND S 18 INVCI n18_CDNS_672673910984 $T=6615 -12785 1 180 $X=5775 $Y=-14805
X27 VDD 7 VDD 10 p18_CDNS_672673910983 $T=-875 -9780 0 0 $X=-1785 $Y=-10210
X28 VDD 12 VDD A p18_CDNS_672673910983 $T=2255 -19050 1 0 $X=1345 $Y=-21280
X29 VDD 12 14 9 p18_CDNS_672673910983 $T=3695 -19050 1 0 $X=2785 $Y=-21280
X30 VDD VDD 17 14 p18_CDNS_672673910983 $T=5635 -19050 1 0 $X=4725 $Y=-21280
X31 VDD VDD 18 11 p18_CDNS_672673910983 $T=5675 -9780 0 0 $X=4765 $Y=-10210
X32 VDD VDD A 21 p18_CDNS_672673910981 $T=-115 -19050 1 0 $X=-1025 $Y=-21280
X33 VDD 11 B 22 p18_CDNS_672673910981 $T=3305 -9780 0 0 $X=2395 $Y=-10210
X34 VDD 9 B 21 p18_CDNS_672673910982 $T=315 -19050 1 0 $X=-240 $Y=-21280
X35 VDD VDD A 22 p18_CDNS_672673910982 $T=3735 -9780 0 0 $X=3180 $Y=-10210
.ENDS
***************************************

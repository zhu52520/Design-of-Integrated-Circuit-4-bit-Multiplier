* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_672340308762 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_672340308760 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT HA_2_3 C A INVC B GND VDD S
** N=11 EP=7 IP=23 FDC=14
M0 GND INVC C GND NM L=1.8e-07 W=2.2e-07 $X=45525 $Y=-24530 $D=0
M1 10 A GND GND NM L=1.8e-07 W=4.4e-07 $X=46285 $Y=-24650 $D=0
M2 INVC B 10 GND NM L=1.8e-07 W=4.4e-07 $X=46715 $Y=-24650 $D=0
M3 GND A 6 GND NM L=1.8e-07 W=4.4e-07 $X=49375 $Y=-24650 $D=0
M4 S 4 GND GND NM L=1.8e-07 W=2.2e-07 $X=52075 $Y=-24640 $D=0
M5 INVC A VDD VDD PM L=1.8e-07 W=4.4e-07 $X=46285 $Y=-21205 $D=4
M6 4 INVC VDD VDD PM L=1.8e-07 W=4.4e-07 $X=48945 $Y=-21205 $D=4
M7 11 A 4 VDD PM L=1.8e-07 W=8.8e-07 $X=49705 $Y=-21645 $D=4
M8 VDD B 11 VDD PM L=1.8e-07 W=8.8e-07 $X=50135 $Y=-21645 $D=4
X9 VDD C VDD INVC p18_CDNS_672340308762 $T=45565 -21205 0 0 $X=44655 $Y=-21635
X10 VDD INVC VDD B p18_CDNS_672340308762 $T=47005 -21205 0 0 $X=46095 $Y=-21635
X11 VDD VDD S 4 p18_CDNS_672340308762 $T=52075 -21205 0 0 $X=51165 $Y=-21635
X12 GND 4 6 INVC n18_CDNS_672340308760 $T=48655 -24650 0 0 $X=47995 $Y=-26670
X13 GND GND 6 B n18_CDNS_672340308760 $T=50095 -24650 0 0 $X=49435 $Y=-26670
.ENDS
***************************************

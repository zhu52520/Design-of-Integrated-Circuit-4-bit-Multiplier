* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673695010463 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673695010462 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673695010460 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT MUX2_SC GND VDD I0 I1 S OUT
** N=12 EP=6 IP=29 FDC=14
M0 OUT 1 4 GND NM L=1.8e-07 W=4.4e-07 $X=-6405 $Y=-10725 $D=0
M1 GND 3 4 GND NM L=1.8e-07 W=4.4e-07 $X=-3745 $Y=-10725 $D=0
M2 11 S VDD VDD PM L=1.8e-07 W=8.8e-07 $X=-7125 $Y=-5465 $D=4
M3 OUT 1 11 VDD PM L=1.8e-07 W=8.8e-07 $X=-6695 $Y=-5465 $D=4
M4 12 2 OUT VDD PM L=1.8e-07 W=8.8e-07 $X=-5975 $Y=-5465 $D=4
M5 VDD 3 12 VDD PM L=1.8e-07 W=8.8e-07 $X=-5545 $Y=-5465 $D=4
X6 VDD 1 I0 p18_CDNS_673695010463 $T=-13145 -5025 0 0 $X=-14055 $Y=-5455
X7 VDD 2 I1 p18_CDNS_673695010463 $T=-11125 -5025 0 0 $X=-12035 $Y=-5455
X8 VDD 3 S p18_CDNS_673695010463 $T=-9105 -5025 0 0 $X=-10015 $Y=-5455
X9 GND 1 I0 n18_CDNS_673695010462 $T=-13145 -10625 0 0 $X=-13845 $Y=-11855
X10 GND 2 I1 n18_CDNS_673695010462 $T=-11125 -10625 0 0 $X=-11825 $Y=-11855
X11 GND 3 S n18_CDNS_673695010462 $T=-9105 -10625 0 0 $X=-9805 $Y=-11855
X12 GND OUT 4 S n18_CDNS_673695010460 $T=-7125 -10725 0 0 $X=-7785 $Y=-11855
X13 GND GND 4 2 n18_CDNS_673695010460 $T=-4465 -10725 0 0 $X=-5125 $Y=-11855
.ENDS
***************************************

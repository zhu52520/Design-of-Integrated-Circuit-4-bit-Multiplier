* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_672672265856 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672672265857 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 3 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_6726722658510 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=6 EP=5 IP=8 FDC=2
X0 1 2 4 6 p18_CDNS_672672265857 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 6 p18_CDNS_6726722658510 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_672672265850 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672672265859 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672672265858 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6
** N=7 EP=6 IP=15 FDC=4
X0 1 5 7 n18_CDNS_672672265850 $T=0 0 0 0 $X=-660 $Y=-2020
X1 1 2 6 7 n18_CDNS_672672265859 $T=430 0 0 0 $X=110 $Y=-2020
X2 1 3 4 2 n18_CDNS_672672265858 $T=2370 0 0 0 $X=1710 $Y=-2020
X3 1 1 4 6 n18_CDNS_672672265858 $T=3810 0 0 0 $X=3150 $Y=-2020
.ENDS
***************************************
.SUBCKT p18_CDNS_672672265852 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_6726722658511 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 3 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672672265851 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_672672265854 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_672672265855 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 3 6 n18_CDNS_672672265855 $T=0 -1580 1 0 $X=-700 $Y=-2150
X1 1 4 5 6 n18_CDNS_672672265855 $T=0 0 0 0 $X=-700 $Y=-1180
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=4
X0 1 1 2 1 3 8 ICV_3 $T=0 0 0 0 $X=-700 $Y=-2150
X1 1 4 6 5 7 8 ICV_3 $T=2020 0 0 0 $X=1320 $Y=-2150
.ENDS
***************************************
.SUBCKT p18_CDNS_672672265853 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT Multiplier X3 O6 Y0 Y1 Y2 Y3 O5 O4 O7 X2 X1 X0 O0 O3 O2 GND VDD O1
** N=187 EP=18 IP=521 FDC=444
M0 GND 5 2 GND NM L=1.8e-07 W=2.2e-07 $X=-1090 $Y=-4200 $D=0
M1 GND 56 3 GND NM L=1.8e-07 W=2.2e-07 $X=-1090 $Y=-480 $D=0
M2 5 7 O7 GND NM L=1.8e-07 W=4.4e-07 $X=-330 $Y=-13550 $D=0
M3 GND 52 35 GND NM L=1.8e-07 W=2.2e-07 $X=1770 $Y=6545 $D=0
M4 GND 53 27 GND NM L=1.8e-07 W=2.2e-07 $X=1770 $Y=8345 $D=0
M5 GND 54 4 GND NM L=1.8e-07 W=2.2e-07 $X=1770 $Y=13165 $D=0
M6 GND 55 8 GND NM L=1.8e-07 W=2.2e-07 $X=1770 $Y=14965 $D=0
M7 GND 3 62 GND NM L=1.8e-07 W=4.4e-07 $X=2760 $Y=-4300 $D=0
M8 GND 4 63 GND NM L=1.8e-07 W=4.4e-07 $X=2760 $Y=-600 $D=0
M9 65 22 7 GND NM L=1.8e-07 W=4.4e-07 $X=3440 $Y=-17250 $D=0
M10 GND 57 65 GND NM L=1.8e-07 W=4.4e-07 $X=4160 $Y=-17250 $D=0
M11 GND 58 64 GND NM L=1.8e-07 W=4.4e-07 $X=4360 $Y=-13550 $D=0
M12 57 11 GND GND NM L=1.8e-07 W=2.2e-07 $X=4920 $Y=-17150 $D=0
M13 155 9 GND GND NM L=1.8e-07 W=4.4e-07 $X=5080 $Y=-13550 $D=0
M14 9 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=5460 $Y=-4200 $D=0
M15 14 60 GND GND NM L=1.8e-07 W=2.2e-07 $X=5460 $Y=-480 $D=0
M16 58 11 155 GND NM L=1.8e-07 W=4.4e-07 $X=5510 $Y=-13550 $D=0
M17 GND 66 46 GND NM L=1.8e-07 W=2.2e-07 $X=6620 $Y=6545 $D=0
M18 GND 67 38 GND NM L=1.8e-07 W=2.2e-07 $X=6620 $Y=8345 $D=0
M19 GND 68 26 GND NM L=1.8e-07 W=2.2e-07 $X=6620 $Y=13165 $D=0
M20 GND 69 10 GND NM L=1.8e-07 W=2.2e-07 $X=6620 $Y=14965 $D=0
M21 GND 87 12 GND NM L=1.8e-07 W=4.4e-07 $X=7440 $Y=-600 $D=0
M22 73 58 71 GND NM L=1.8e-07 W=4.4e-07 $X=7450 $Y=-13550 $D=0
M23 GND 74 11 GND NM L=1.8e-07 W=2.2e-07 $X=7480 $Y=-4200 $D=0
M24 156 11 79 GND NM L=1.8e-07 W=4.4e-07 $X=7700 $Y=-17250 $D=0
M25 GND 9 156 GND NM L=1.8e-07 W=4.4e-07 $X=8130 $Y=-17250 $D=0
M26 GND 9 73 GND NM L=1.8e-07 W=4.4e-07 $X=8170 $Y=-13550 $D=0
M27 79 57 GND GND NM L=1.8e-07 W=2.2e-07 $X=8890 $Y=-17150 $D=0
M28 73 11 GND GND NM L=1.8e-07 W=4.4e-07 $X=8890 $Y=-13550 $D=0
M29 GND 27 83 GND NM L=1.8e-07 W=4.4e-07 $X=9380 $Y=-600 $D=0
M30 157 27 GND GND NM L=1.8e-07 W=4.4e-07 $X=10100 $Y=-600 $D=0
M31 87 26 157 GND NM L=1.8e-07 W=4.4e-07 $X=10530 $Y=-600 $D=0
M32 80 79 GND GND NM L=1.8e-07 W=4.4e-07 $X=10870 $Y=-17250 $D=0
M33 81 71 GND GND NM L=1.8e-07 W=4.4e-07 $X=10870 $Y=-13550 $D=0
M34 83 21 87 GND NM L=1.8e-07 W=4.4e-07 $X=11250 $Y=-600 $D=0
M35 GND 12 85 GND NM L=1.8e-07 W=4.4e-07 $X=11330 $Y=-4300 $D=0
M36 GND 75 49 GND NM L=1.8e-07 W=2.2e-07 $X=11470 $Y=6545 $D=0
M37 GND 76 13 GND NM L=1.8e-07 W=2.2e-07 $X=11470 $Y=8345 $D=0
M38 GND 77 24 GND NM L=1.8e-07 W=2.2e-07 $X=11470 $Y=13165 $D=0
M39 GND 78 21 GND NM L=1.8e-07 W=2.2e-07 $X=11470 $Y=14965 $D=0
M40 O6 22 80 GND NM L=1.8e-07 W=4.4e-07 $X=11630 $Y=-17250 $D=0
M41 GND 26 83 GND NM L=1.8e-07 W=4.4e-07 $X=11970 $Y=-600 $D=0
M42 158 26 GND GND NM L=1.8e-07 W=4.4e-07 $X=12690 $Y=-600 $D=0
M43 159 27 158 GND NM L=1.8e-07 W=4.4e-07 $X=13120 $Y=-600 $D=0
M44 99 21 159 GND NM L=1.8e-07 W=4.4e-07 $X=13550 $Y=-600 $D=0
M45 25 82 GND GND NM L=1.8e-07 W=2.2e-07 $X=14030 $Y=-4200 $D=0
M46 96 87 99 GND NM L=1.8e-07 W=4.4e-07 $X=14270 $Y=-600 $D=0
M47 GND 21 96 GND NM L=1.8e-07 W=4.4e-07 $X=14990 $Y=-600 $D=0
M48 98 34 22 GND NM L=1.8e-07 W=4.4e-07 $X=15510 $Y=-17250 $D=0
M49 96 27 GND GND NM L=1.8e-07 W=4.4e-07 $X=15710 $Y=-600 $D=0
M50 GND 107 28 GND NM L=1.8e-07 W=4.4e-07 $X=16010 $Y=-4300 $D=0
M51 GND 92 98 GND NM L=1.8e-07 W=4.4e-07 $X=16230 $Y=-17250 $D=0
M52 GND 88 O0 GND NM L=1.8e-07 W=2.2e-07 $X=16320 $Y=6545 $D=0
M53 GND 89 50 GND NM L=1.8e-07 W=2.2e-07 $X=16320 $Y=8345 $D=0
M54 GND 90 45 GND NM L=1.8e-07 W=2.2e-07 $X=16320 $Y=13165 $D=0
M55 GND 91 23 GND NM L=1.8e-07 W=2.2e-07 $X=16320 $Y=14965 $D=0
M56 GND 93 95 GND NM L=1.8e-07 W=4.4e-07 $X=16430 $Y=-13550 $D=0
M57 GND 26 96 GND NM L=1.8e-07 W=4.4e-07 $X=16430 $Y=-600 $D=0
M58 92 28 GND GND NM L=1.8e-07 W=2.2e-07 $X=16990 $Y=-17150 $D=0
M59 160 25 GND GND NM L=1.8e-07 W=4.4e-07 $X=17150 $Y=-13550 $D=0
M60 29 99 GND GND NM L=1.8e-07 W=4.4e-07 $X=17150 $Y=-600 $D=0
M61 93 28 160 GND NM L=1.8e-07 W=4.4e-07 $X=17580 $Y=-13550 $D=0
M62 GND 31 101 GND NM L=1.8e-07 W=4.4e-07 $X=17950 $Y=-4300 $D=0
M63 161 31 GND GND NM L=1.8e-07 W=4.4e-07 $X=18670 $Y=-4300 $D=0
M64 107 33 161 GND NM L=1.8e-07 W=4.4e-07 $X=19100 $Y=-4300 $D=0
M65 GND 104 33 GND NM L=1.8e-07 W=2.2e-07 $X=19130 $Y=-480 $D=0
M66 105 93 102 GND NM L=1.8e-07 W=4.4e-07 $X=19520 $Y=-13550 $D=0
M67 162 28 106 GND NM L=1.8e-07 W=4.4e-07 $X=19770 $Y=-17250 $D=0
M68 101 29 107 GND NM L=1.8e-07 W=4.4e-07 $X=19820 $Y=-4300 $D=0
M69 GND 25 162 GND NM L=1.8e-07 W=4.4e-07 $X=20200 $Y=-17250 $D=0
M70 GND 25 105 GND NM L=1.8e-07 W=4.4e-07 $X=20240 $Y=-13550 $D=0
M71 GND 33 101 GND NM L=1.8e-07 W=4.4e-07 $X=20540 $Y=-4300 $D=0
M72 106 92 GND GND NM L=1.8e-07 W=2.2e-07 $X=20960 $Y=-17150 $D=0
M73 105 28 GND GND NM L=1.8e-07 W=4.4e-07 $X=20960 $Y=-13550 $D=0
M74 163 33 GND GND NM L=1.8e-07 W=4.4e-07 $X=21260 $Y=-4300 $D=0
M75 164 31 163 GND NM L=1.8e-07 W=4.4e-07 $X=21690 $Y=-4300 $D=0
M76 114 29 164 GND NM L=1.8e-07 W=4.4e-07 $X=22120 $Y=-4300 $D=0
M77 113 107 114 GND NM L=1.8e-07 W=4.4e-07 $X=22840 $Y=-4300 $D=0
M78 109 106 GND GND NM L=1.8e-07 W=4.4e-07 $X=22940 $Y=-17250 $D=0
M79 110 102 GND GND NM L=1.8e-07 W=4.4e-07 $X=22940 $Y=-13550 $D=0
M80 GND 24 111 GND NM L=1.8e-07 W=4.4e-07 $X=22980 $Y=-600 $D=0
M81 GND 29 113 GND NM L=1.8e-07 W=4.4e-07 $X=23560 $Y=-4300 $D=0
M82 O5 34 109 GND NM L=1.8e-07 W=4.4e-07 $X=23700 $Y=-17250 $D=0
M83 113 31 GND GND NM L=1.8e-07 W=4.4e-07 $X=24280 $Y=-4300 $D=0
M84 GND 33 113 GND NM L=1.8e-07 W=4.4e-07 $X=25000 $Y=-4300 $D=0
M85 42 108 GND GND NM L=1.8e-07 W=2.2e-07 $X=25680 $Y=-480 $D=0
M86 36 114 GND GND NM L=1.8e-07 W=4.4e-07 $X=25720 $Y=-4300 $D=0
M87 120 118 34 GND NM L=1.8e-07 W=4.4e-07 $X=27580 $Y=-17250 $D=0
M88 GND 130 37 GND NM L=1.8e-07 W=4.4e-07 $X=27660 $Y=-4300 $D=0
M89 GND 121 31 GND NM L=1.8e-07 W=2.2e-07 $X=27700 $Y=-480 $D=0
M90 GND 115 120 GND NM L=1.8e-07 W=4.4e-07 $X=28300 $Y=-17250 $D=0
M91 GND 116 119 GND NM L=1.8e-07 W=4.4e-07 $X=28500 $Y=-13550 $D=0
M92 115 37 GND GND NM L=1.8e-07 W=2.2e-07 $X=29060 $Y=-17150 $D=0
M93 165 36 GND GND NM L=1.8e-07 W=4.4e-07 $X=29220 $Y=-13550 $D=0
M94 GND 40 124 GND NM L=1.8e-07 W=4.4e-07 $X=29600 $Y=-4300 $D=0
M95 116 37 165 GND NM L=1.8e-07 W=4.4e-07 $X=29650 $Y=-13550 $D=0
M96 166 40 GND GND NM L=1.8e-07 W=4.4e-07 $X=30320 $Y=-4300 $D=0
M97 130 42 166 GND NM L=1.8e-07 W=4.4e-07 $X=30750 $Y=-4300 $D=0
M98 124 39 130 GND NM L=1.8e-07 W=4.4e-07 $X=31470 $Y=-4300 $D=0
M99 GND 35 126 GND NM L=1.8e-07 W=4.4e-07 $X=31550 $Y=-600 $D=0
M100 128 116 125 GND NM L=1.8e-07 W=4.4e-07 $X=31590 $Y=-13550 $D=0
M101 167 37 129 GND NM L=1.8e-07 W=4.4e-07 $X=31840 $Y=-17250 $D=0
M102 GND 42 124 GND NM L=1.8e-07 W=4.4e-07 $X=32190 $Y=-4300 $D=0
M103 GND 36 167 GND NM L=1.8e-07 W=4.4e-07 $X=32270 $Y=-17250 $D=0
M104 GND 36 128 GND NM L=1.8e-07 W=4.4e-07 $X=32310 $Y=-13550 $D=0
M105 168 42 GND GND NM L=1.8e-07 W=4.4e-07 $X=32910 $Y=-4300 $D=0
M106 129 115 GND GND NM L=1.8e-07 W=2.2e-07 $X=33030 $Y=-17150 $D=0
M107 128 37 GND GND NM L=1.8e-07 W=4.4e-07 $X=33030 $Y=-13550 $D=0
M108 169 40 168 GND NM L=1.8e-07 W=4.4e-07 $X=33340 $Y=-4300 $D=0
M109 135 39 169 GND NM L=1.8e-07 W=4.4e-07 $X=33770 $Y=-4300 $D=0
M110 40 122 GND GND NM L=1.8e-07 W=2.2e-07 $X=34250 $Y=-480 $D=0
M111 134 130 135 GND NM L=1.8e-07 W=4.4e-07 $X=34490 $Y=-4300 $D=0
M112 131 129 GND GND NM L=1.8e-07 W=4.4e-07 $X=35010 $Y=-17250 $D=0
M113 132 125 GND GND NM L=1.8e-07 W=4.4e-07 $X=35010 $Y=-13550 $D=0
M114 GND 39 134 GND NM L=1.8e-07 W=4.4e-07 $X=35210 $Y=-4300 $D=0
M115 O4 118 131 GND NM L=1.8e-07 W=4.4e-07 $X=35770 $Y=-17250 $D=0
M116 134 40 GND GND NM L=1.8e-07 W=4.4e-07 $X=35930 $Y=-4300 $D=0
M117 GND 141 39 GND NM L=1.8e-07 W=4.4e-07 $X=36230 $Y=-600 $D=0
M118 GND 42 134 GND NM L=1.8e-07 W=4.4e-07 $X=36650 $Y=-4300 $D=0
M119 44 135 GND GND NM L=1.8e-07 W=4.4e-07 $X=37370 $Y=-4300 $D=0
M120 GND 117 118 GND NM L=1.8e-07 W=2.2e-07 $X=37750 $Y=-13430 $D=0
M121 GND 46 136 GND NM L=1.8e-07 W=4.4e-07 $X=38170 $Y=-600 $D=0
M122 170 46 GND GND NM L=1.8e-07 W=4.4e-07 $X=38890 $Y=-600 $D=0
M123 141 13 170 GND NM L=1.8e-07 W=4.4e-07 $X=39320 $Y=-600 $D=0
M124 GND 138 43 GND NM L=1.8e-07 W=2.2e-07 $X=39350 $Y=-4200 $D=0
M125 136 45 141 GND NM L=1.8e-07 W=4.4e-07 $X=40040 $Y=-600 $D=0
M126 GND 13 136 GND NM L=1.8e-07 W=4.4e-07 $X=40760 $Y=-600 $D=0
M127 171 13 GND GND NM L=1.8e-07 W=4.4e-07 $X=41480 $Y=-600 $D=0
M128 GND 43 140 GND NM L=1.8e-07 W=4.4e-07 $X=41600 $Y=-13550 $D=0
M129 172 46 171 GND NM L=1.8e-07 W=4.4e-07 $X=41910 $Y=-600 $D=0
M130 147 45 172 GND NM L=1.8e-07 W=4.4e-07 $X=42340 $Y=-600 $D=0
M131 145 141 147 GND NM L=1.8e-07 W=4.4e-07 $X=43060 $Y=-600 $D=0
M132 GND 48 143 GND NM L=1.8e-07 W=4.4e-07 $X=43200 $Y=-4300 $D=0
M133 GND 45 145 GND NM L=1.8e-07 W=4.4e-07 $X=43780 $Y=-600 $D=0
M134 O3 139 GND GND NM L=1.8e-07 W=2.2e-07 $X=44300 $Y=-13430 $D=0
M135 145 46 GND GND NM L=1.8e-07 W=4.4e-07 $X=44500 $Y=-600 $D=0
M136 GND 13 145 GND NM L=1.8e-07 W=4.4e-07 $X=45220 $Y=-600 $D=0
M137 O2 142 GND GND NM L=1.8e-07 W=2.2e-07 $X=45900 $Y=-4200 $D=0
M138 47 147 GND GND NM L=1.8e-07 W=4.4e-07 $X=45940 $Y=-600 $D=0
M139 GND 149 48 GND NM L=1.8e-07 W=2.2e-07 $X=47920 $Y=-480 $D=0
M140 GND 49 151 GND NM L=1.8e-07 W=4.4e-07 $X=51770 $Y=-600 $D=0
M141 O1 150 GND GND NM L=1.8e-07 W=2.2e-07 $X=54470 $Y=-480 $D=0
M142 5 6 O7 VDD PM L=1.8e-07 W=4.4e-07 $X=-330 $Y=-10105 $D=4
M143 5 3 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-330 $Y=-7745 $D=4
M144 56 4 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-330 $Y=2845 $D=4
M145 35 52 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=970 $Y=5205 $D=4
M146 GND X3 35 VDD PM L=1.8e-07 W=2.2e-07 $X=1770 $Y=5205 $D=4
M147 GND X3 27 VDD PM L=1.8e-07 W=2.2e-07 $X=1770 $Y=9685 $D=4
M148 GND X3 4 VDD PM L=1.8e-07 W=2.2e-07 $X=1770 $Y=11825 $D=4
M149 GND X3 8 VDD PM L=1.8e-07 W=2.2e-07 $X=1770 $Y=16305 $D=4
M150 59 5 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=2330 $Y=-7745 $D=4
M151 60 56 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=2330 $Y=2845 $D=4
M152 VDD 8 173 VDD PM L=1.8e-07 W=8.8e-07 $X=3520 $Y=-7745 $D=4
M153 64 22 7 VDD PM L=1.8e-07 W=4.4e-07 $X=3560 $Y=-10105 $D=4
M154 66 X2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=3800 $Y=5085 $D=4
M155 VDD 57 65 VDD PM L=1.8e-07 W=8.8e-07 $X=4360 $Y=-20695 $D=4
M156 58 9 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=5080 $Y=-10105 $D=4
M157 VDD 11 58 VDD PM L=1.8e-07 W=4.4e-07 $X=5800 $Y=-10105 $D=4
M158 46 66 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=5820 $Y=5205 $D=4
M159 GND X2 46 VDD PM L=1.8e-07 W=2.2e-07 $X=6620 $Y=5205 $D=4
M160 GND X2 38 VDD PM L=1.8e-07 W=2.2e-07 $X=6620 $Y=9685 $D=4
M161 GND X2 26 VDD PM L=1.8e-07 W=2.2e-07 $X=6620 $Y=11825 $D=4
M162 GND X2 10 VDD PM L=1.8e-07 W=2.2e-07 $X=6620 $Y=16305 $D=4
M163 VDD 87 12 VDD PM L=1.8e-07 W=8.8e-07 $X=7440 $Y=2405 $D=4
M164 71 58 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=7740 $Y=-10105 $D=4
M165 72 9 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=8170 $Y=-20695 $D=4
M166 74 12 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=8240 $Y=-7745 $D=4
M167 VDD 11 174 VDD PM L=1.8e-07 W=8.8e-07 $X=8930 $Y=-10545 $D=4
M168 VDD 14 74 VDD PM L=1.8e-07 W=4.4e-07 $X=8960 $Y=-7745 $D=4
M169 VDD 27 84 VDD PM L=1.8e-07 W=8.8e-07 $X=9380 $Y=2405 $D=4
M170 175 27 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10100 $Y=2405 $D=4
M171 87 26 175 VDD PM L=1.8e-07 W=8.8e-07 $X=10530 $Y=2405 $D=4
M172 81 71 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=10870 $Y=-10545 $D=4
M173 82 74 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=10900 $Y=-7745 $D=4
M174 84 21 87 VDD PM L=1.8e-07 W=8.8e-07 $X=11250 $Y=2405 $D=4
M175 GND X1 49 VDD PM L=1.8e-07 W=2.2e-07 $X=11470 $Y=5205 $D=4
M176 GND X1 13 VDD PM L=1.8e-07 W=2.2e-07 $X=11470 $Y=9685 $D=4
M177 GND X1 24 VDD PM L=1.8e-07 W=2.2e-07 $X=11470 $Y=11825 $D=4
M178 GND X1 21 VDD PM L=1.8e-07 W=2.2e-07 $X=11470 $Y=16305 $D=4
M179 O6 16 80 VDD PM L=1.8e-07 W=4.4e-07 $X=11590 $Y=-20695 $D=4
M180 O6 22 81 VDD PM L=1.8e-07 W=4.4e-07 $X=11630 $Y=-10105 $D=4
M181 VDD 26 84 VDD PM L=1.8e-07 W=8.8e-07 $X=11970 $Y=2405 $D=4
M182 VDD 14 176 VDD PM L=1.8e-07 W=8.8e-07 $X=12090 $Y=-7745 $D=4
M183 177 26 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=12690 $Y=2405 $D=4
M184 178 27 177 VDD PM L=1.8e-07 W=8.8e-07 $X=13120 $Y=2405 $D=4
M185 99 21 178 VDD PM L=1.8e-07 W=8.8e-07 $X=13550 $Y=2405 $D=4
M186 93 34 16 VDD PM L=1.8e-07 W=4.4e-07 $X=13680 $Y=-10105 $D=4
M187 97 87 99 VDD PM L=1.8e-07 W=8.8e-07 $X=14270 $Y=2405 $D=4
M188 VDD 21 97 VDD PM L=1.8e-07 W=8.8e-07 $X=14990 $Y=2405 $D=4
M189 95 34 22 VDD PM L=1.8e-07 W=4.4e-07 $X=15630 $Y=-10105 $D=4
M190 97 27 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=15710 $Y=2405 $D=4
M191 VDD 107 28 VDD PM L=1.8e-07 W=8.8e-07 $X=16010 $Y=-7745 $D=4
M192 GND X0 O0 VDD PM L=1.8e-07 W=2.2e-07 $X=16320 $Y=5205 $D=4
M193 GND X0 50 VDD PM L=1.8e-07 W=2.2e-07 $X=16320 $Y=9685 $D=4
M194 GND X0 45 VDD PM L=1.8e-07 W=2.2e-07 $X=16320 $Y=11825 $D=4
M195 GND X0 23 VDD PM L=1.8e-07 W=2.2e-07 $X=16320 $Y=16305 $D=4
M196 VDD 92 98 VDD PM L=1.8e-07 W=8.8e-07 $X=16430 $Y=-20695 $D=4
M197 VDD 26 97 VDD PM L=1.8e-07 W=8.8e-07 $X=16430 $Y=2405 $D=4
M198 93 25 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=17150 $Y=-10105 $D=4
M199 29 99 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=17150 $Y=2405 $D=4
M200 VDD 31 100 VDD PM L=1.8e-07 W=8.8e-07 $X=17950 $Y=-7745 $D=4
M201 179 31 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=18670 $Y=-7745 $D=4
M202 107 33 179 VDD PM L=1.8e-07 W=8.8e-07 $X=19100 $Y=-7745 $D=4
M203 102 93 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=19810 $Y=-10105 $D=4
M204 100 29 107 VDD PM L=1.8e-07 W=8.8e-07 $X=19820 $Y=-7745 $D=4
M205 104 24 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=19890 $Y=2845 $D=4
M206 103 25 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=20240 $Y=-20695 $D=4
M207 VDD 33 100 VDD PM L=1.8e-07 W=8.8e-07 $X=20540 $Y=-7745 $D=4
M208 180 33 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=21260 $Y=-7745 $D=4
M209 181 31 180 VDD PM L=1.8e-07 W=8.8e-07 $X=21690 $Y=-7745 $D=4
M210 114 29 181 VDD PM L=1.8e-07 W=8.8e-07 $X=22120 $Y=-7745 $D=4
M211 108 104 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=22550 $Y=2845 $D=4
M212 112 107 114 VDD PM L=1.8e-07 W=8.8e-07 $X=22840 $Y=-7745 $D=4
M213 110 102 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=22940 $Y=-10545 $D=4
M214 VDD 29 112 VDD PM L=1.8e-07 W=8.8e-07 $X=23560 $Y=-7745 $D=4
M215 O5 32 109 VDD PM L=1.8e-07 W=4.4e-07 $X=23660 $Y=-20695 $D=4
M216 O5 34 110 VDD PM L=1.8e-07 W=4.4e-07 $X=23700 $Y=-10105 $D=4
M217 112 31 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=24280 $Y=-7745 $D=4
M218 VDD 33 112 VDD PM L=1.8e-07 W=8.8e-07 $X=25000 $Y=-7745 $D=4
M219 36 114 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=25720 $Y=-7745 $D=4
M220 VDD 130 37 VDD PM L=1.8e-07 W=8.8e-07 $X=27660 $Y=-7745 $D=4
M221 119 118 34 VDD PM L=1.8e-07 W=4.4e-07 $X=27700 $Y=-10105 $D=4
M222 121 35 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=28460 $Y=2845 $D=4
M223 VDD 115 120 VDD PM L=1.8e-07 W=8.8e-07 $X=28500 $Y=-20695 $D=4
M224 116 36 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=29220 $Y=-10105 $D=4
M225 VDD 40 123 VDD PM L=1.8e-07 W=8.8e-07 $X=29600 $Y=-7745 $D=4
M226 182 40 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=30320 $Y=-7745 $D=4
M227 130 42 182 VDD PM L=1.8e-07 W=8.8e-07 $X=30750 $Y=-7745 $D=4
M228 122 121 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31120 $Y=2845 $D=4
M229 123 39 130 VDD PM L=1.8e-07 W=8.8e-07 $X=31470 $Y=-7745 $D=4
M230 125 116 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31880 $Y=-10105 $D=4
M231 VDD 42 123 VDD PM L=1.8e-07 W=8.8e-07 $X=32190 $Y=-7745 $D=4
M232 127 36 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=32310 $Y=-20695 $D=4
M233 183 42 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=32910 $Y=-7745 $D=4
M234 184 40 183 VDD PM L=1.8e-07 W=8.8e-07 $X=33340 $Y=-7745 $D=4
M235 135 39 184 VDD PM L=1.8e-07 W=8.8e-07 $X=33770 $Y=-7745 $D=4
M236 133 130 135 VDD PM L=1.8e-07 W=8.8e-07 $X=34490 $Y=-7745 $D=4
M237 VDD 39 133 VDD PM L=1.8e-07 W=8.8e-07 $X=35210 $Y=-7745 $D=4
M238 O4 117 131 VDD PM L=1.8e-07 W=4.4e-07 $X=35730 $Y=-20695 $D=4
M239 O4 118 132 VDD PM L=1.8e-07 W=4.4e-07 $X=35770 $Y=-10105 $D=4
M240 133 40 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35930 $Y=-7745 $D=4
M241 VDD 141 39 VDD PM L=1.8e-07 W=8.8e-07 $X=36230 $Y=2405 $D=4
M242 VDD 42 133 VDD PM L=1.8e-07 W=8.8e-07 $X=36650 $Y=-7745 $D=4
M243 44 135 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=37370 $Y=-7745 $D=4
M244 VDD 46 137 VDD PM L=1.8e-07 W=8.8e-07 $X=38170 $Y=2405 $D=4
M245 117 43 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=38510 $Y=-10105 $D=4
M246 185 46 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=38890 $Y=2405 $D=4
M247 VDD 44 117 VDD PM L=1.8e-07 W=4.4e-07 $X=39230 $Y=-10105 $D=4
M248 141 13 185 VDD PM L=1.8e-07 W=8.8e-07 $X=39320 $Y=2405 $D=4
M249 137 45 141 VDD PM L=1.8e-07 W=8.8e-07 $X=40040 $Y=2405 $D=4
M250 138 48 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=40110 $Y=-7745 $D=4
M251 VDD 13 137 VDD PM L=1.8e-07 W=8.8e-07 $X=40760 $Y=2405 $D=4
M252 139 117 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=41170 $Y=-10105 $D=4
M253 186 13 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41480 $Y=2405 $D=4
M254 187 46 186 VDD PM L=1.8e-07 W=8.8e-07 $X=41910 $Y=2405 $D=4
M255 147 45 187 VDD PM L=1.8e-07 W=8.8e-07 $X=42340 $Y=2405 $D=4
M256 142 138 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=42770 $Y=-7745 $D=4
M257 146 141 147 VDD PM L=1.8e-07 W=8.8e-07 $X=43060 $Y=2405 $D=4
M258 VDD 45 146 VDD PM L=1.8e-07 W=8.8e-07 $X=43780 $Y=2405 $D=4
M259 O3 139 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=44300 $Y=-10105 $D=4
M260 146 46 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44500 $Y=2405 $D=4
M261 VDD 13 146 VDD PM L=1.8e-07 W=8.8e-07 $X=45220 $Y=2405 $D=4
M262 47 147 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=45940 $Y=2405 $D=4
M263 149 49 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=48680 $Y=2845 $D=4
M264 150 149 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=51340 $Y=2845 $D=4
X265 VDD 2 O7 7 p18_CDNS_672672265856 $T=-1050 -10105 0 0 $X=-1960 $Y=-10535
X266 VDD 2 VDD 5 p18_CDNS_672672265856 $T=-1050 -7305 1 0 $X=-1960 $Y=-9095
X267 VDD 3 VDD 56 p18_CDNS_672672265856 $T=-1050 2845 0 0 $X=-1960 $Y=2415
X268 VDD 5 VDD 8 p18_CDNS_672672265856 $T=390 -7305 1 0 $X=-520 $Y=-9095
X269 VDD 56 VDD 10 p18_CDNS_672672265856 $T=390 2845 0 0 $X=-520 $Y=2415
X270 VDD 6 58 22 p18_CDNS_672672265856 $T=1610 -10105 0 0 $X=700 $Y=-10535
X271 VDD 57 6 16 p18_CDNS_672672265856 $T=1840 -20255 0 180 $X=750 $Y=-22045
X272 VDD 65 7 16 p18_CDNS_672672265856 $T=3780 -20255 0 180 $X=2690 $Y=-22045
X273 VDD VDD 9 59 p18_CDNS_672672265856 $T=5460 -7305 1 0 $X=4550 $Y=-9095
X274 VDD VDD 14 60 p18_CDNS_672672265856 $T=5460 2845 0 0 $X=4550 $Y=2415
X275 VDD 11 VDD 74 p18_CDNS_672672265856 $T=7520 -7305 1 0 $X=6610 $Y=-9095
X276 VDD 92 16 32 p18_CDNS_672672265856 $T=13910 -20255 0 180 $X=12820 $Y=-22045
X277 VDD VDD 25 82 p18_CDNS_672672265856 $T=14030 -7305 1 0 $X=13120 $Y=-9095
X278 VDD 98 22 32 p18_CDNS_672672265856 $T=15850 -20255 0 180 $X=14760 $Y=-22045
X279 VDD 93 VDD 28 p18_CDNS_672672265856 $T=17870 -10105 0 0 $X=16960 $Y=-10535
X280 VDD 33 VDD 104 p18_CDNS_672672265856 $T=19170 2845 0 0 $X=18260 $Y=2415
X281 VDD 104 VDD 23 p18_CDNS_672672265856 $T=20610 2845 0 0 $X=19700 $Y=2415
X282 VDD VDD 42 108 p18_CDNS_672672265856 $T=25680 2845 0 0 $X=24770 $Y=2415
X283 VDD 32 116 118 p18_CDNS_672672265856 $T=25750 -10105 0 0 $X=24840 $Y=-10535
X284 VDD 115 32 117 p18_CDNS_672672265856 $T=25980 -20255 0 180 $X=24890 $Y=-22045
X285 VDD 120 34 117 p18_CDNS_672672265856 $T=27920 -20255 0 180 $X=26830 $Y=-22045
X286 VDD 31 VDD 121 p18_CDNS_672672265856 $T=27740 2845 0 0 $X=26830 $Y=2415
X287 VDD 121 VDD 38 p18_CDNS_672672265856 $T=29180 2845 0 0 $X=28270 $Y=2415
X288 VDD 116 VDD 37 p18_CDNS_672672265856 $T=29940 -10105 0 0 $X=29030 $Y=-10535
X289 VDD VDD 40 122 p18_CDNS_672672265856 $T=34250 2845 0 0 $X=33340 $Y=2415
X290 VDD 118 VDD 117 p18_CDNS_672672265856 $T=37790 -10105 0 0 $X=36880 $Y=-10535
X291 VDD 43 VDD 138 p18_CDNS_672672265856 $T=39390 -7305 1 0 $X=38480 $Y=-9095
X292 VDD 138 VDD 47 p18_CDNS_672672265856 $T=40830 -7305 1 0 $X=39920 $Y=-9095
X293 VDD VDD O2 142 p18_CDNS_672672265856 $T=45900 -7305 1 0 $X=44990 $Y=-9095
X294 VDD 48 VDD 149 p18_CDNS_672672265856 $T=47960 2845 0 0 $X=47050 $Y=2415
X295 VDD 149 VDD 50 p18_CDNS_672672265856 $T=49400 2845 0 0 $X=48490 $Y=2415
X296 VDD VDD O1 150 p18_CDNS_672672265856 $T=54470 2845 0 0 $X=53560 $Y=2415
X297 VDD 59 3 173 p18_CDNS_672672265857 $T=3090 -6865 1 0 $X=2180 $Y=-9095
X298 VDD 71 9 174 p18_CDNS_672672265857 $T=8500 -10545 0 0 $X=7590 $Y=-10975
X299 VDD 82 12 176 p18_CDNS_672672265857 $T=11660 -6865 1 0 $X=10750 $Y=-9095
X300 VDD 60 VDD 4 10 ICV_1 $T=3090 2405 0 0 $X=2180 $Y=1975
X301 VDD VDD 57 11 9 ICV_1 $T=5080 -19815 1 0 $X=4170 $Y=-22045
X302 VDD VDD 92 28 25 ICV_1 $T=17150 -19815 1 0 $X=16240 $Y=-22045
X303 VDD 102 VDD 25 28 ICV_1 $T=20570 -10545 0 0 $X=19660 $Y=-10975
X304 VDD 108 VDD 24 23 ICV_1 $T=23310 2405 0 0 $X=22400 $Y=1975
X305 VDD VDD 115 37 36 ICV_1 $T=29220 -19815 1 0 $X=28310 $Y=-22045
X306 VDD 122 VDD 35 38 ICV_1 $T=31880 2405 0 0 $X=30970 $Y=1975
X307 VDD 125 VDD 36 37 ICV_1 $T=32640 -10545 0 0 $X=31730 $Y=-10975
X308 VDD 139 VDD 43 44 ICV_1 $T=41930 -10545 0 0 $X=41020 $Y=-10975
X309 VDD 142 VDD 48 47 ICV_1 $T=43530 -6865 1 0 $X=42620 $Y=-9095
X310 VDD 150 VDD 49 50 ICV_1 $T=52100 2405 0 0 $X=51190 $Y=1975
X311 GND 2 O7 6 n18_CDNS_672672265858 $T=-1050 -13550 0 0 $X=-1710 $Y=-15570
X312 GND 58 6 16 n18_CDNS_672672265858 $T=1790 -13550 1 180 $X=950 $Y=-15570
X313 GND 64 7 16 n18_CDNS_672672265858 $T=3740 -13550 1 180 $X=2900 $Y=-15570
X314 GND O6 81 16 n18_CDNS_672672265858 $T=11810 -13550 1 180 $X=10970 $Y=-15570
X315 GND 93 16 32 n18_CDNS_672672265858 $T=13860 -13550 1 180 $X=13020 $Y=-15570
X316 GND 95 22 32 n18_CDNS_672672265858 $T=15810 -13550 1 180 $X=14970 $Y=-15570
X317 GND O5 110 32 n18_CDNS_672672265858 $T=23880 -13550 1 180 $X=23040 $Y=-15570
X318 GND 116 32 117 n18_CDNS_672672265858 $T=25930 -13550 1 180 $X=25090 $Y=-15570
X319 GND 119 34 117 n18_CDNS_672672265858 $T=27880 -13550 1 180 $X=27040 $Y=-15570
X320 GND O4 132 117 n18_CDNS_672672265858 $T=35950 -13550 1 180 $X=35110 $Y=-15570
X321 GND 5 59 62 3 8 ICV_2 $T=-330 -3860 1 0 $X=-990 $Y=-4650
X322 GND 56 60 63 4 10 ICV_2 $T=-330 -600 0 0 $X=-990 $Y=-2620
X323 GND 74 82 85 12 14 ICV_2 $T=8240 -3860 1 0 $X=7580 $Y=-4650
X324 GND 104 108 111 24 23 ICV_2 $T=19890 -600 0 0 $X=19230 $Y=-2620
X325 GND 121 122 126 35 38 ICV_2 $T=28460 -600 0 0 $X=27800 $Y=-2620
X326 GND 117 139 140 43 44 ICV_2 $T=38510 -13550 0 0 $X=37850 $Y=-15570
X327 GND 138 142 143 48 47 ICV_2 $T=40110 -3860 1 0 $X=39450 $Y=-4650
X328 GND 149 150 151 49 50 ICV_2 $T=48680 -600 0 0 $X=48020 $Y=-2620
X329 VDD 64 VDD 58 p18_CDNS_672672265852 $T=4320 -10545 0 0 $X=3410 $Y=-10975
X330 VDD 72 VDD 11 p18_CDNS_672672265852 $T=7450 -19815 1 0 $X=6540 $Y=-22045
X331 VDD 72 79 57 p18_CDNS_672672265852 $T=8890 -19815 1 0 $X=7980 $Y=-22045
X332 VDD VDD 80 79 p18_CDNS_672672265852 $T=10830 -19815 1 0 $X=9920 $Y=-22045
X333 VDD 95 VDD 93 p18_CDNS_672672265852 $T=16390 -10545 0 0 $X=15480 $Y=-10975
X334 VDD 103 VDD 28 p18_CDNS_672672265852 $T=19520 -19815 1 0 $X=18610 $Y=-22045
X335 VDD 103 106 92 p18_CDNS_672672265852 $T=20960 -19815 1 0 $X=20050 $Y=-22045
X336 VDD VDD 109 106 p18_CDNS_672672265852 $T=22900 -19815 1 0 $X=21990 $Y=-22045
X337 VDD 119 VDD 116 p18_CDNS_672672265852 $T=28460 -10545 0 0 $X=27550 $Y=-10975
X338 VDD 127 VDD 37 p18_CDNS_672672265852 $T=31590 -19815 1 0 $X=30680 $Y=-22045
X339 VDD 127 129 115 p18_CDNS_672672265852 $T=33030 -19815 1 0 $X=32120 $Y=-22045
X340 VDD VDD 131 129 p18_CDNS_672672265852 $T=34970 -19815 1 0 $X=34060 $Y=-22045
X341 VDD VDD 132 125 p18_CDNS_672672265852 $T=35010 -10545 0 0 $X=34100 $Y=-10975
X342 GND 57 9 n18_CDNS_6726722658511 $T=5720 -16930 1 0 $X=5020 $Y=-17500
X343 GND 92 25 n18_CDNS_6726722658511 $T=17790 -16930 1 0 $X=17090 $Y=-17500
X344 GND 115 36 n18_CDNS_6726722658511 $T=29860 -16930 1 0 $X=29160 $Y=-17500
X345 6 57 22 GND n18_CDNS_672672265851 $T=1500 -16810 1 0 $X=840 $Y=-17600
X346 16 92 34 GND n18_CDNS_672672265851 $T=13570 -16810 1 0 $X=12910 $Y=-17600
X347 32 115 118 GND n18_CDNS_672672265851 $T=25640 -16810 1 0 $X=24980 $Y=-17600
X348 VDD Y1 27 53 p18_CDNS_672672265854 $T=970 9685 0 0 $X=20 $Y=9155
X349 VDD Y2 4 54 p18_CDNS_672672265854 $T=970 12045 1 0 $X=20 $Y=10475
X350 VDD Y3 8 55 p18_CDNS_672672265854 $T=970 16305 0 0 $X=20 $Y=15775
X351 VDD Y1 38 67 p18_CDNS_672672265854 $T=5820 9685 0 0 $X=4870 $Y=9155
X352 VDD Y2 26 68 p18_CDNS_672672265854 $T=5820 12045 1 0 $X=4870 $Y=10475
X353 VDD Y3 10 69 p18_CDNS_672672265854 $T=5820 16305 0 0 $X=4870 $Y=15775
X354 VDD Y0 49 75 p18_CDNS_672672265854 $T=10670 5425 1 0 $X=9720 $Y=3855
X355 VDD Y1 13 76 p18_CDNS_672672265854 $T=10670 9685 0 0 $X=9720 $Y=9155
X356 VDD Y2 24 77 p18_CDNS_672672265854 $T=10670 12045 1 0 $X=9720 $Y=10475
X357 VDD Y3 21 78 p18_CDNS_672672265854 $T=10670 16305 0 0 $X=9720 $Y=15775
X358 VDD Y0 O0 88 p18_CDNS_672672265854 $T=15520 5425 1 0 $X=14570 $Y=3855
X359 VDD Y1 50 89 p18_CDNS_672672265854 $T=15520 9685 0 0 $X=14570 $Y=9155
X360 VDD Y2 45 90 p18_CDNS_672672265854 $T=15520 12045 1 0 $X=14570 $Y=10475
X361 VDD Y3 23 91 p18_CDNS_672672265854 $T=15520 16305 0 0 $X=14570 $Y=15775
X362 GND 53 52 Y1 Y0 27 35 X3 ICV_4 $T=-1050 6765 1 0 $X=-1750 $Y=6195
X363 GND 55 54 Y3 Y2 8 4 X3 ICV_4 $T=-1050 13385 1 0 $X=-1750 $Y=12815
X364 GND 67 66 Y1 Y0 38 46 X2 ICV_4 $T=3800 6765 1 0 $X=3100 $Y=6195
X365 GND 69 68 Y3 Y2 10 26 X2 ICV_4 $T=3800 13385 1 0 $X=3100 $Y=12815
X366 GND 76 75 Y1 Y0 13 49 X1 ICV_4 $T=8650 6765 1 0 $X=7950 $Y=6195
X367 GND 78 77 Y3 Y2 21 24 X1 ICV_4 $T=8650 13385 1 0 $X=7950 $Y=12815
X368 GND 89 88 Y1 Y0 50 O0 X0 ICV_4 $T=13500 6765 1 0 $X=12800 $Y=6195
X369 GND 91 90 Y3 Y2 23 45 X0 ICV_4 $T=13500 13385 1 0 $X=12800 $Y=12815
X370 VDD 52 X3 p18_CDNS_672672265853 $T=-1050 5525 1 0 $X=-1960 $Y=3855
X371 VDD 53 X3 p18_CDNS_672672265853 $T=-1050 9585 0 0 $X=-1960 $Y=9155
X372 VDD 54 X3 p18_CDNS_672672265853 $T=-1050 12145 1 0 $X=-1960 $Y=10475
X373 VDD 55 X3 p18_CDNS_672672265853 $T=-1050 16205 0 0 $X=-1960 $Y=15775
X374 VDD 67 X2 p18_CDNS_672672265853 $T=3800 9585 0 0 $X=2890 $Y=9155
X375 VDD 68 X2 p18_CDNS_672672265853 $T=3800 12145 1 0 $X=2890 $Y=10475
X376 VDD 69 X2 p18_CDNS_672672265853 $T=3800 16205 0 0 $X=2890 $Y=15775
X377 VDD 75 X1 p18_CDNS_672672265853 $T=8650 5525 1 0 $X=7740 $Y=3855
X378 VDD 76 X1 p18_CDNS_672672265853 $T=8650 9585 0 0 $X=7740 $Y=9155
X379 VDD 77 X1 p18_CDNS_672672265853 $T=8650 12145 1 0 $X=7740 $Y=10475
X380 VDD 78 X1 p18_CDNS_672672265853 $T=8650 16205 0 0 $X=7740 $Y=15775
X381 VDD 88 X0 p18_CDNS_672672265853 $T=13500 5525 1 0 $X=12590 $Y=3855
X382 VDD 89 X0 p18_CDNS_672672265853 $T=13500 9585 0 0 $X=12590 $Y=9155
X383 VDD 90 X0 p18_CDNS_672672265853 $T=13500 12145 1 0 $X=12590 $Y=10475
X384 VDD 91 X0 p18_CDNS_672672265853 $T=13500 16205 0 0 $X=12590 $Y=15775
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_672748097267 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 1 3 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672748097262 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672748097263 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 4 2 3 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_672748097261 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=8 EP=5 IP=14 FDC=3
X0 1 3 7 p18_CDNS_672748097262 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 7 8 p18_CDNS_672748097263 $T=430 0 0 0 $X=-125 $Y=-430
X2 1 2 5 8 p18_CDNS_672748097261 $T=860 0 0 0 $X=305 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_672748097264 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 3 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672748097265 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_672748097266 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 3 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=8 EP=7 IP=15 FDC=4
X0 1 1 2 8 n18_CDNS_672748097264 $T=0 0 0 0 $X=-660 $Y=-1350
X1 1 2 5 7 n18_CDNS_672748097264 $T=2370 0 0 0 $X=1710 $Y=-1350
X2 1 3 5 8 n18_CDNS_672748097265 $T=430 0 0 0 $X=110 $Y=-1350
X3 1 4 6 n18_CDNS_672748097266 $T=4240 0 0 0 $X=3580 $Y=-1350
.ENDS
***************************************
.SUBCKT p18_CDNS_672748097260 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT Register_9bit INVQ0 CLK Q0 RST D0 INVQ1 Q1 D1 INVQ2 Q2 D2 INVQ3 Q3 D3 INVQ4 Q4 D4 INVQ5 Q5 D5
+ INVQ6 Q6 D6 INVQ7 Q7 D7 INVQ8 Q8 D8 VDD GND
** N=67 EP=31 IP=189 FDC=135
M0 GND Q0 INVQ0 GND NM L=1.8e-07 W=4.4e-07 $X=-63620 $Y=-10560 $D=0
M1 GND 5 59 GND NM L=1.8e-07 W=4.4e-07 $X=-60100 $Y=-10560 $D=0
M2 5 7 GND GND NM L=1.8e-07 W=4.4e-07 $X=-59380 $Y=-10560 $D=0
M3 GND D0 7 GND NM L=1.8e-07 W=2.2e-07 $X=-56680 $Y=-10440 $D=0
M4 GND Q1 INVQ1 GND NM L=1.8e-07 W=4.4e-07 $X=-54700 $Y=-10560 $D=0
M5 GND 12 60 GND NM L=1.8e-07 W=4.4e-07 $X=-51180 $Y=-10560 $D=0
M6 12 13 GND GND NM L=1.8e-07 W=4.4e-07 $X=-50460 $Y=-10560 $D=0
M7 GND D1 13 GND NM L=1.8e-07 W=2.2e-07 $X=-47760 $Y=-10440 $D=0
M8 GND Q2 INVQ2 GND NM L=1.8e-07 W=4.4e-07 $X=-45780 $Y=-10560 $D=0
M9 GND 18 61 GND NM L=1.8e-07 W=4.4e-07 $X=-42260 $Y=-10560 $D=0
M10 18 19 GND GND NM L=1.8e-07 W=4.4e-07 $X=-41540 $Y=-10560 $D=0
M11 GND D2 19 GND NM L=1.8e-07 W=2.2e-07 $X=-38840 $Y=-10440 $D=0
M12 GND Q3 INVQ3 GND NM L=1.8e-07 W=4.4e-07 $X=-36860 $Y=-10560 $D=0
M13 GND 24 62 GND NM L=1.8e-07 W=4.4e-07 $X=-33340 $Y=-10560 $D=0
M14 24 25 GND GND NM L=1.8e-07 W=4.4e-07 $X=-32620 $Y=-10560 $D=0
M15 GND D3 25 GND NM L=1.8e-07 W=2.2e-07 $X=-29920 $Y=-10440 $D=0
M16 GND Q4 INVQ4 GND NM L=1.8e-07 W=4.4e-07 $X=-27940 $Y=-10560 $D=0
M17 GND 30 63 GND NM L=1.8e-07 W=4.4e-07 $X=-24420 $Y=-10560 $D=0
M18 30 31 GND GND NM L=1.8e-07 W=4.4e-07 $X=-23700 $Y=-10560 $D=0
M19 GND D4 31 GND NM L=1.8e-07 W=2.2e-07 $X=-21000 $Y=-10440 $D=0
M20 GND Q5 INVQ5 GND NM L=1.8e-07 W=4.4e-07 $X=-19020 $Y=-10560 $D=0
M21 GND 36 64 GND NM L=1.8e-07 W=4.4e-07 $X=-15500 $Y=-10560 $D=0
M22 36 37 GND GND NM L=1.8e-07 W=4.4e-07 $X=-14780 $Y=-10560 $D=0
M23 GND D5 37 GND NM L=1.8e-07 W=2.2e-07 $X=-12080 $Y=-10440 $D=0
M24 GND Q6 INVQ6 GND NM L=1.8e-07 W=4.4e-07 $X=-10100 $Y=-10560 $D=0
M25 GND 42 65 GND NM L=1.8e-07 W=4.4e-07 $X=-6580 $Y=-10560 $D=0
M26 42 43 GND GND NM L=1.8e-07 W=4.4e-07 $X=-5860 $Y=-10560 $D=0
M27 GND D6 43 GND NM L=1.8e-07 W=2.2e-07 $X=-3160 $Y=-10440 $D=0
M28 GND Q7 INVQ7 GND NM L=1.8e-07 W=4.4e-07 $X=-1180 $Y=-10560 $D=0
M29 GND 48 66 GND NM L=1.8e-07 W=4.4e-07 $X=2340 $Y=-10560 $D=0
M30 48 49 GND GND NM L=1.8e-07 W=4.4e-07 $X=3060 $Y=-10560 $D=0
M31 GND D7 49 GND NM L=1.8e-07 W=2.2e-07 $X=5760 $Y=-10440 $D=0
M32 GND Q8 INVQ8 GND NM L=1.8e-07 W=4.4e-07 $X=7740 $Y=-10560 $D=0
M33 GND 54 67 GND NM L=1.8e-07 W=4.4e-07 $X=11260 $Y=-10560 $D=0
M34 54 55 GND GND NM L=1.8e-07 W=4.4e-07 $X=11980 $Y=-10560 $D=0
M35 GND D8 55 GND NM L=1.8e-07 W=2.2e-07 $X=14680 $Y=-10440 $D=0
M36 VDD Q0 INVQ0 VDD PM L=1.8e-07 W=8.8e-07 $X=-63620 $Y=-8480 $D=4
M37 VDD CLK 4 VDD PM L=1.8e-07 W=8.8e-07 $X=-60200 $Y=-8480 $D=4
M38 VDD Q1 INVQ1 VDD PM L=1.8e-07 W=8.8e-07 $X=-54700 $Y=-8480 $D=4
M39 VDD CLK 11 VDD PM L=1.8e-07 W=8.8e-07 $X=-51280 $Y=-8480 $D=4
M40 VDD Q2 INVQ2 VDD PM L=1.8e-07 W=8.8e-07 $X=-45780 $Y=-8480 $D=4
M41 VDD CLK 17 VDD PM L=1.8e-07 W=8.8e-07 $X=-42360 $Y=-8480 $D=4
M42 VDD Q3 INVQ3 VDD PM L=1.8e-07 W=8.8e-07 $X=-36860 $Y=-8480 $D=4
M43 VDD CLK 23 VDD PM L=1.8e-07 W=8.8e-07 $X=-33440 $Y=-8480 $D=4
M44 VDD Q4 INVQ4 VDD PM L=1.8e-07 W=8.8e-07 $X=-27940 $Y=-8480 $D=4
M45 VDD CLK 29 VDD PM L=1.8e-07 W=8.8e-07 $X=-24520 $Y=-8480 $D=4
M46 VDD Q5 INVQ5 VDD PM L=1.8e-07 W=8.8e-07 $X=-19020 $Y=-8480 $D=4
M47 VDD CLK 35 VDD PM L=1.8e-07 W=8.8e-07 $X=-15600 $Y=-8480 $D=4
M48 VDD Q6 INVQ6 VDD PM L=1.8e-07 W=8.8e-07 $X=-10100 $Y=-8480 $D=4
M49 VDD CLK 41 VDD PM L=1.8e-07 W=8.8e-07 $X=-6680 $Y=-8480 $D=4
M50 VDD Q7 INVQ7 VDD PM L=1.8e-07 W=8.8e-07 $X=-1180 $Y=-8480 $D=4
M51 VDD CLK 47 VDD PM L=1.8e-07 W=8.8e-07 $X=2240 $Y=-8480 $D=4
M52 VDD Q8 INVQ8 VDD PM L=1.8e-07 W=8.8e-07 $X=7740 $Y=-8480 $D=4
M53 VDD CLK 53 VDD PM L=1.8e-07 W=8.8e-07 $X=11160 $Y=-8480 $D=4
X54 VDD 7 D0 p18_CDNS_672748097267 $T=-56680 -8040 0 0 $X=-57590 $Y=-8470
X55 VDD 13 D1 p18_CDNS_672748097267 $T=-47760 -8040 0 0 $X=-48670 $Y=-8470
X56 VDD 19 D2 p18_CDNS_672748097267 $T=-38840 -8040 0 0 $X=-39750 $Y=-8470
X57 VDD 25 D3 p18_CDNS_672748097267 $T=-29920 -8040 0 0 $X=-30830 $Y=-8470
X58 VDD 31 D4 p18_CDNS_672748097267 $T=-21000 -8040 0 0 $X=-21910 $Y=-8470
X59 VDD 37 D5 p18_CDNS_672748097267 $T=-12080 -8040 0 0 $X=-12990 $Y=-8470
X60 VDD 43 D6 p18_CDNS_672748097267 $T=-3160 -8040 0 0 $X=-4070 $Y=-8470
X61 VDD 49 D7 p18_CDNS_672748097267 $T=5760 -8040 0 0 $X=4850 $Y=-8470
X62 VDD 55 D8 p18_CDNS_672748097267 $T=14680 -8040 0 0 $X=13770 $Y=-8470
X63 VDD 5 7 RST CLK ICV_1 $T=-59480 -8480 0 0 $X=-60390 $Y=-8910
X64 VDD 12 13 RST CLK ICV_1 $T=-50560 -8480 0 0 $X=-51470 $Y=-8910
X65 VDD 18 19 RST CLK ICV_1 $T=-41640 -8480 0 0 $X=-42550 $Y=-8910
X66 VDD 24 25 RST CLK ICV_1 $T=-32720 -8480 0 0 $X=-33630 $Y=-8910
X67 VDD 30 31 RST CLK ICV_1 $T=-23800 -8480 0 0 $X=-24710 $Y=-8910
X68 VDD 36 37 RST CLK ICV_1 $T=-14880 -8480 0 0 $X=-15790 $Y=-8910
X69 VDD 42 43 RST CLK ICV_1 $T=-5960 -8480 0 0 $X=-6870 $Y=-8910
X70 VDD 48 49 RST CLK ICV_1 $T=2960 -8480 0 0 $X=2050 $Y=-8910
X71 VDD 54 55 RST CLK ICV_1 $T=11880 -8480 0 0 $X=10970 $Y=-8910
X72 GND 4 Q0 5 CLK RST 59 ICV_2 $T=-62900 -10560 0 0 $X=-63560 $Y=-11910
X73 GND 11 Q1 12 CLK RST 60 ICV_2 $T=-53980 -10560 0 0 $X=-54640 $Y=-11910
X74 GND 17 Q2 18 CLK RST 61 ICV_2 $T=-45060 -10560 0 0 $X=-45720 $Y=-11910
X75 GND 23 Q3 24 CLK RST 62 ICV_2 $T=-36140 -10560 0 0 $X=-36800 $Y=-11910
X76 GND 29 Q4 30 CLK RST 63 ICV_2 $T=-27220 -10560 0 0 $X=-27880 $Y=-11910
X77 GND 35 Q5 36 CLK RST 64 ICV_2 $T=-18300 -10560 0 0 $X=-18960 $Y=-11910
X78 GND 41 Q6 42 CLK RST 65 ICV_2 $T=-9380 -10560 0 0 $X=-10040 $Y=-11910
X79 GND 47 Q7 48 CLK RST 66 ICV_2 $T=-460 -10560 0 0 $X=-1120 $Y=-11910
X80 GND 53 Q8 54 CLK RST 67 ICV_2 $T=8460 -10560 0 0 $X=7800 $Y=-11910
X81 VDD Q0 4 p18_CDNS_672748097260 $T=-62900 -8480 0 0 $X=-63810 $Y=-8910
X82 VDD Q1 11 p18_CDNS_672748097260 $T=-53980 -8480 0 0 $X=-54890 $Y=-8910
X83 VDD Q2 17 p18_CDNS_672748097260 $T=-45060 -8480 0 0 $X=-45970 $Y=-8910
X84 VDD Q3 23 p18_CDNS_672748097260 $T=-36140 -8480 0 0 $X=-37050 $Y=-8910
X85 VDD Q4 29 p18_CDNS_672748097260 $T=-27220 -8480 0 0 $X=-28130 $Y=-8910
X86 VDD Q5 35 p18_CDNS_672748097260 $T=-18300 -8480 0 0 $X=-19210 $Y=-8910
X87 VDD Q6 41 p18_CDNS_672748097260 $T=-9380 -8480 0 0 $X=-10290 $Y=-8910
X88 VDD Q7 47 p18_CDNS_672748097260 $T=-460 -8480 0 0 $X=-1370 $Y=-8910
X89 VDD Q8 53 p18_CDNS_672748097260 $T=8460 -8480 0 0 $X=7550 $Y=-8910
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT TSPC_v2 CLK Q RST D VDD GND
** N=13 EP=6 IP=0 FDC=13
M0 10 3 GND GND NM L=1.8e-07 W=4.4e-07 $X=40330 $Y=-13745 $D=0
M1 Q CLK 10 GND NM L=1.8e-07 W=4.4e-07 $X=40760 $Y=-13745 $D=0
M2 11 CLK 3 GND NM L=1.8e-07 W=4.4e-07 $X=42700 $Y=-13745 $D=0
M3 GND 4 11 GND NM L=1.8e-07 W=4.4e-07 $X=43130 $Y=-13745 $D=0
M4 4 6 GND GND NM L=1.8e-07 W=4.4e-07 $X=43850 $Y=-13745 $D=0
M5 GND RST 4 GND NM L=1.8e-07 W=4.4e-07 $X=44570 $Y=-13745 $D=0
M6 GND D 6 GND NM L=1.8e-07 W=2.2e-07 $X=46550 $Y=-13625 $D=0
M7 Q 3 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=40330 $Y=-10740 $D=4
M8 VDD CLK 3 VDD PM L=1.8e-07 W=8.8e-07 $X=43030 $Y=-10740 $D=4
M9 12 6 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=43750 $Y=-10740 $D=4
M10 13 RST 12 VDD PM L=1.8e-07 W=8.8e-07 $X=44180 $Y=-10740 $D=4
M11 4 CLK 13 VDD PM L=1.8e-07 W=8.8e-07 $X=44610 $Y=-10740 $D=4
M12 VDD D 6 VDD PM L=1.8e-07 W=4.4e-07 $X=46550 $Y=-10300 $D=4
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673696248871 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT n18_CDNS_673696248870 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Buffer2 GND VDD X Y
** N=5 EP=4 IP=14 FDC=4
X0 VDD 4 X p18_CDNS_673696248871 $T=42130 -20700 0 0 $X=41220 $Y=-21130
X1 VDD Y 4 p18_CDNS_673696248871 $T=44150 -20700 0 0 $X=43240 $Y=-21130
X2 GND 4 X n18_CDNS_673696248870 $T=42130 -26300 0 0 $X=41430 $Y=-27530
X3 GND Y 4 n18_CDNS_673696248870 $T=44150 -26300 0 0 $X=43450 $Y=-27530
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673547882912 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT Bitcell BIT INVBIT GND WL VDD
** N=7 EP=5 IP=10 FDC=6
M0 4 6 GND GND NM L=1.8e-07 W=8e-07 $X=25290 $Y=-15850 $D=0
M1 4 WL BIT GND NM L=1.8e-07 W=4.4e-07 $X=25340 $Y=-17480 $D=0
M2 6 WL INVBIT GND NM L=1.8e-07 W=4.4e-07 $X=27000 $Y=-17480 $D=0
M3 GND 4 6 GND NM L=1.8e-07 W=8e-07 $X=27310 $Y=-15850 $D=0
X4 VDD VDD 4 6 p18_CDNS_673547882912 $T=25290 -13900 0 0 $X=24340 $Y=-14430
X5 VDD 6 VDD 4 p18_CDNS_673547882912 $T=27310 -13900 0 0 $X=26360 $Y=-14430
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT p18_CDNS_673868691721 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673868691723 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 4 3 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673868691728 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=6 EP=5 IP=8 FDC=2
X0 1 2 4 6 p18_CDNS_673868691723 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 5 6 p18_CDNS_673868691728 $T=430 0 0 0 $X=-125 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_673868691722 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 3 2 1 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673868691727 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 4 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673868691726 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6
** N=7 EP=6 IP=15 FDC=4
X0 1 5 7 n18_CDNS_673868691722 $T=0 0 0 0 $X=-660 $Y=-2020
X1 1 2 6 7 n18_CDNS_673868691727 $T=430 0 0 0 $X=110 $Y=-2020
X2 1 3 4 2 n18_CDNS_673868691726 $T=2370 0 0 0 $X=1710 $Y=-2020
X3 1 1 4 6 n18_CDNS_673868691726 $T=3810 0 0 0 $X=3150 $Y=-2020
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4
** N=4 EP=4 IP=8 FDC=2
X0 1 2 1 3 p18_CDNS_673868691721 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 1 4 p18_CDNS_673868691721 $T=1440 0 0 0 $X=530 $Y=-430
.ENDS
***************************************
.SUBCKT p18_CDNS_6738686917210 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=8.8e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=2
X0 1 2 1 4 p18_CDNS_6738686917210 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 2 3 5 p18_CDNS_6738686917210 $T=1440 0 0 0 $X=530 $Y=-430
.ENDS
***************************************
.SUBCKT n18_CDNS_6738686917211 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 1 3 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673868691729 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 NM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 3 6 n18_CDNS_673868691726 $T=-1950 0 0 0 $X=-2610 $Y=-2020
X1 1 4 5 6 n18_CDNS_673868691726 $T=0 0 0 0 $X=-660 $Y=-2020
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=3
X0 1 2 3 7 n18_CDNS_673868691726 $T=0 0 0 0 $X=-660 $Y=-2020
X1 1 4 5 6 7 8 ICV_5 $T=-2050 0 0 0 $X=-4660 $Y=-2020
.ENDS
***************************************
.SUBCKT n18_CDNS_673868691725 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6
** N=6 EP=6 IP=8 FDC=2
X0 1 2 3 6 n18_CDNS_673868691725 $T=0 -1580 1 0 $X=-700 $Y=-2150
X1 1 4 5 6 n18_CDNS_673868691725 $T=0 0 0 0 $X=-700 $Y=-1180
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=4
X0 1 1 2 1 3 8 ICV_7 $T=0 0 0 0 $X=-700 $Y=-2150
X1 1 4 6 5 7 8 ICV_7 $T=2020 0 0 0 $X=1320 $Y=-2150
.ENDS
***************************************
.SUBCKT p18_CDNS_673868691720 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673868691724 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 PM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=4
X0 1 2 8 p18_CDNS_673868691720 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 8 p18_CDNS_673868691720 $T=0 2560 1 0 $X=-910 $Y=890
X2 1 4 5 2 p18_CDNS_673868691724 $T=2020 100 0 0 $X=1070 $Y=-430
X3 1 6 7 3 p18_CDNS_673868691724 $T=2020 2460 1 0 $X=1070 $Y=890
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5
** N=5 EP=5 IP=7 FDC=2
X0 1 2 5 p18_CDNS_673868691720 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 3 4 2 p18_CDNS_673868691724 $T=2020 100 0 0 $X=1070 $Y=-430
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=4
X0 1 2 3 4 7 ICV_10 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 5 3 6 8 ICV_10 $T=4850 0 0 0 $X=3940 $Y=-430
.ENDS
***************************************
.SUBCKT VU_reg Q8I Q7I Q6I Q3I Q5I Q2I Q4I Q1I Q0I B3 X3 A3 A2 A1 A0 Y0 Y1 Y2 Y3 RST
+ CLK B2 X2 B1 X1 B0 X0 Q3 Q8 INVQ3 INVQ8 Q2 Q7 INVQ2 INVQ7 Q1 Q6 INVQ1 INVQ6 Q0
+ Q5 INVQ0 INVQ5 Q4 INVQ4 GND VDD
** N=572 EP=47 IP=1168 FDC=1313
M0 135 37 Q8I GND NM L=1.8e-07 W=4.4e-07 $X=30420 $Y=-20465 $D=0
M1 GND 144 14 GND NM L=1.8e-07 W=2.2e-07 $X=30500 $Y=-46265 $D=0
M2 GND 18 12 GND NM L=1.8e-07 W=2.2e-07 $X=30500 $Y=-42545 $D=0
M3 GND 19 13 GND NM L=1.8e-07 W=2.2e-07 $X=30500 $Y=5535 $D=0
M4 GND 145 15 GND NM L=1.8e-07 W=2.2e-07 $X=30500 $Y=9255 $D=0
M5 GND 146 135 GND NM L=1.8e-07 W=4.4e-07 $X=31140 $Y=-20465 $D=0
M6 18 23 27 GND NM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-33415 $D=0
M7 19 24 20 GND NM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-3815 $D=0
M8 GND 147 134 GND NM L=1.8e-07 W=4.4e-07 $X=31340 $Y=-16765 $D=0
M9 146 27 GND GND NM L=1.8e-07 W=2.2e-07 $X=31900 $Y=-20365 $D=0
M10 449 20 GND GND NM L=1.8e-07 W=4.4e-07 $X=32060 $Y=-16765 $D=0
M11 147 27 449 GND NM L=1.8e-07 W=4.4e-07 $X=32490 $Y=-16765 $D=0
M12 GND 136 25 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-61710 $D=0
M13 GND 137 16 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-59910 $D=0
M14 GND 138 66 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-55090 $D=0
M15 GND 139 83 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-53290 $D=0
M16 GND 140 85 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=16280 $D=0
M17 GND 141 67 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=18080 $D=0
M18 GND 142 17 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=22900 $D=0
M19 GND 143 26 GND NM L=1.8e-07 W=2.2e-07 $X=33360 $Y=24700 $D=0
M20 GND 16 159 GND NM L=1.8e-07 W=4.4e-07 $X=34350 $Y=-46365 $D=0
M21 GND 14 160 GND NM L=1.8e-07 W=4.4e-07 $X=34350 $Y=-42665 $D=0
M22 GND 15 161 GND NM L=1.8e-07 W=4.4e-07 $X=34350 $Y=5435 $D=0
M23 GND 17 162 GND NM L=1.8e-07 W=4.4e-07 $X=34350 $Y=9135 $D=0
M24 176 147 158 GND NM L=1.8e-07 W=4.4e-07 $X=34430 $Y=-16765 $D=0
M25 450 27 177 GND NM L=1.8e-07 W=4.4e-07 $X=34680 $Y=-20465 $D=0
M26 166 55 23 GND NM L=1.8e-07 W=4.4e-07 $X=35030 $Y=-29715 $D=0
M27 167 56 24 GND NM L=1.8e-07 W=4.4e-07 $X=35030 $Y=-7515 $D=0
M28 GND 20 450 GND NM L=1.8e-07 W=4.4e-07 $X=35110 $Y=-20465 $D=0
M29 GND 20 176 GND NM L=1.8e-07 W=4.4e-07 $X=35150 $Y=-16765 $D=0
M30 GND 148 166 GND NM L=1.8e-07 W=4.4e-07 $X=35750 $Y=-29715 $D=0
M31 GND 149 167 GND NM L=1.8e-07 W=4.4e-07 $X=35750 $Y=-7515 $D=0
M32 177 146 GND GND NM L=1.8e-07 W=2.2e-07 $X=35870 $Y=-20365 $D=0
M33 176 27 GND GND NM L=1.8e-07 W=4.4e-07 $X=35870 $Y=-16765 $D=0
M34 GND 150 163 GND NM L=1.8e-07 W=4.4e-07 $X=35950 $Y=-33415 $D=0
M35 GND 151 165 GND NM L=1.8e-07 W=4.4e-07 $X=35950 $Y=-3815 $D=0
M36 148 32 GND GND NM L=1.8e-07 W=2.2e-07 $X=36510 $Y=-29595 $D=0
M37 149 33 GND GND NM L=1.8e-07 W=2.2e-07 $X=36510 $Y=-7415 $D=0
M38 451 28 GND GND NM L=1.8e-07 W=4.4e-07 $X=36670 $Y=-33415 $D=0
M39 452 29 GND GND NM L=1.8e-07 W=4.4e-07 $X=36670 $Y=-3815 $D=0
M40 40 152 GND GND NM L=1.8e-07 W=2.2e-07 $X=37050 $Y=-46265 $D=0
M41 28 153 GND GND NM L=1.8e-07 W=2.2e-07 $X=37050 $Y=-42545 $D=0
M42 29 154 GND GND NM L=1.8e-07 W=2.2e-07 $X=37050 $Y=5535 $D=0
M43 41 155 GND GND NM L=1.8e-07 W=2.2e-07 $X=37050 $Y=9255 $D=0
M44 150 32 451 GND NM L=1.8e-07 W=4.4e-07 $X=37100 $Y=-33415 $D=0
M45 151 33 452 GND NM L=1.8e-07 W=4.4e-07 $X=37100 $Y=-3815 $D=0
M46 178 177 GND GND NM L=1.8e-07 W=4.4e-07 $X=37850 $Y=-20465 $D=0
M47 179 158 GND GND NM L=1.8e-07 W=4.4e-07 $X=37850 $Y=-16765 $D=0
M48 GND 168 30 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-61710 $D=0
M49 GND 169 64 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-59910 $D=0
M50 GND 170 91 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-55090 $D=0
M51 GND 171 108 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-53290 $D=0
M52 GND 172 109 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=16280 $D=0
M53 GND 173 92 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=18080 $D=0
M54 GND 174 65 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=22900 $D=0
M55 GND 175 31 GND NM L=1.8e-07 W=2.2e-07 $X=38210 $Y=24700 $D=0
M56 Q7I 37 178 GND NM L=1.8e-07 W=4.4e-07 $X=38610 $Y=-20465 $D=0
M57 GND 218 34 GND NM L=1.8e-07 W=4.4e-07 $X=39030 $Y=-46365 $D=0
M58 GND 219 35 GND NM L=1.8e-07 W=4.4e-07 $X=39030 $Y=9135 $D=0
M59 186 150 182 GND NM L=1.8e-07 W=4.4e-07 $X=39040 $Y=-33415 $D=0
M60 187 151 183 GND NM L=1.8e-07 W=4.4e-07 $X=39040 $Y=-3815 $D=0
M61 GND 188 32 GND NM L=1.8e-07 W=2.2e-07 $X=39070 $Y=-42545 $D=0
M62 GND 189 33 GND NM L=1.8e-07 W=2.2e-07 $X=39070 $Y=5535 $D=0
M63 453 32 198 GND NM L=1.8e-07 W=4.4e-07 $X=39290 $Y=-29715 $D=0
M64 454 33 199 GND NM L=1.8e-07 W=4.4e-07 $X=39290 $Y=-7515 $D=0
M65 GND 28 453 GND NM L=1.8e-07 W=4.4e-07 $X=39720 $Y=-29715 $D=0
M66 GND 29 454 GND NM L=1.8e-07 W=4.4e-07 $X=39720 $Y=-7515 $D=0
M67 GND 28 186 GND NM L=1.8e-07 W=4.4e-07 $X=39760 $Y=-33415 $D=0
M68 GND 29 187 GND NM L=1.8e-07 W=4.4e-07 $X=39760 $Y=-3815 $D=0
M69 186 32 GND GND NM L=1.8e-07 W=4.4e-07 $X=40480 $Y=-33415 $D=0
M70 198 148 GND GND NM L=1.8e-07 W=2.2e-07 $X=40480 $Y=-29595 $D=0
M71 199 149 GND GND NM L=1.8e-07 W=2.2e-07 $X=40480 $Y=-7415 $D=0
M72 187 33 GND GND NM L=1.8e-07 W=4.4e-07 $X=40480 $Y=-3815 $D=0
M73 GND 66 211 GND NM L=1.8e-07 W=4.4e-07 $X=40970 $Y=-46365 $D=0
M74 GND 67 212 GND NM L=1.8e-07 W=4.4e-07 $X=40970 $Y=9135 $D=0
M75 455 66 GND GND NM L=1.8e-07 W=4.4e-07 $X=41690 $Y=-46365 $D=0
M76 456 67 GND GND NM L=1.8e-07 W=4.4e-07 $X=41690 $Y=9135 $D=0
M77 218 64 455 GND NM L=1.8e-07 W=4.4e-07 $X=42120 $Y=-46365 $D=0
M78 219 65 456 GND NM L=1.8e-07 W=4.4e-07 $X=42120 $Y=9135 $D=0
M79 204 182 GND GND NM L=1.8e-07 W=4.4e-07 $X=42460 $Y=-33415 $D=0
M80 202 198 GND GND NM L=1.8e-07 W=4.4e-07 $X=42460 $Y=-29715 $D=0
M81 203 199 GND GND NM L=1.8e-07 W=4.4e-07 $X=42460 $Y=-7515 $D=0
M82 205 183 GND GND NM L=1.8e-07 W=4.4e-07 $X=42460 $Y=-3815 $D=0
M83 207 71 37 GND NM L=1.8e-07 W=4.4e-07 $X=42490 $Y=-20465 $D=0
M84 211 53 218 GND NM L=1.8e-07 W=4.4e-07 $X=42840 $Y=-46365 $D=0
M85 212 54 219 GND NM L=1.8e-07 W=4.4e-07 $X=42840 $Y=9135 $D=0
M86 GND 34 214 GND NM L=1.8e-07 W=4.4e-07 $X=42920 $Y=-42665 $D=0
M87 GND 35 215 GND NM L=1.8e-07 W=4.4e-07 $X=42920 $Y=5435 $D=0
M88 GND 190 53 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-61710 $D=0
M89 GND 191 60 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-59910 $D=0
M90 GND 192 38 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-55090 $D=0
M91 GND 193 116 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-53290 $D=0
M92 GND 194 117 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=16280 $D=0
M93 GND 195 39 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=18080 $D=0
M94 GND 196 61 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=22900 $D=0
M95 GND 197 54 GND NM L=1.8e-07 W=2.2e-07 $X=43060 $Y=24700 $D=0
M96 GND 200 207 GND NM L=1.8e-07 W=4.4e-07 $X=43210 $Y=-20465 $D=0
M97 59 55 202 GND NM L=1.8e-07 W=4.4e-07 $X=43220 $Y=-29715 $D=0
M98 42 56 203 GND NM L=1.8e-07 W=4.4e-07 $X=43220 $Y=-7515 $D=0
M99 GND 201 206 GND NM L=1.8e-07 W=4.4e-07 $X=43410 $Y=-16765 $D=0
M100 GND 64 211 GND NM L=1.8e-07 W=4.4e-07 $X=43560 $Y=-46365 $D=0
M101 GND 65 212 GND NM L=1.8e-07 W=4.4e-07 $X=43560 $Y=9135 $D=0
M102 200 59 GND GND NM L=1.8e-07 W=2.2e-07 $X=43970 $Y=-20365 $D=0
M103 457 42 GND GND NM L=1.8e-07 W=4.4e-07 $X=44130 $Y=-16765 $D=0
M104 458 64 GND GND NM L=1.8e-07 W=4.4e-07 $X=44280 $Y=-46365 $D=0
M105 459 65 GND GND NM L=1.8e-07 W=4.4e-07 $X=44280 $Y=9135 $D=0
M106 201 59 457 GND NM L=1.8e-07 W=4.4e-07 $X=44560 $Y=-16765 $D=0
M107 460 66 458 GND NM L=1.8e-07 W=4.4e-07 $X=44710 $Y=-46365 $D=0
M108 461 67 459 GND NM L=1.8e-07 W=4.4e-07 $X=44710 $Y=9135 $D=0
M109 243 53 460 GND NM L=1.8e-07 W=4.4e-07 $X=45140 $Y=-46365 $D=0
M110 244 54 461 GND NM L=1.8e-07 W=4.4e-07 $X=45140 $Y=9135 $D=0
M111 62 208 GND GND NM L=1.8e-07 W=2.2e-07 $X=45620 $Y=-42545 $D=0
M112 63 209 GND GND NM L=1.8e-07 W=2.2e-07 $X=45620 $Y=5535 $D=0
M113 237 218 243 GND NM L=1.8e-07 W=4.4e-07 $X=45860 $Y=-46365 $D=0
M114 238 219 244 GND NM L=1.8e-07 W=4.4e-07 $X=45860 $Y=9135 $D=0
M115 242 201 232 GND NM L=1.8e-07 W=4.4e-07 $X=46500 $Y=-16765 $D=0
M116 GND 53 237 GND NM L=1.8e-07 W=4.4e-07 $X=46580 $Y=-46365 $D=0
M117 GND 54 238 GND NM L=1.8e-07 W=4.4e-07 $X=46580 $Y=9135 $D=0
M118 462 59 245 GND NM L=1.8e-07 W=4.4e-07 $X=46750 $Y=-20465 $D=0
M119 240 81 55 GND NM L=1.8e-07 W=4.4e-07 $X=47100 $Y=-29715 $D=0
M120 241 82 56 GND NM L=1.8e-07 W=4.4e-07 $X=47100 $Y=-7515 $D=0
M121 GND 42 462 GND NM L=1.8e-07 W=4.4e-07 $X=47180 $Y=-20465 $D=0
M122 GND 42 242 GND NM L=1.8e-07 W=4.4e-07 $X=47220 $Y=-16765 $D=0
M123 237 66 GND GND NM L=1.8e-07 W=4.4e-07 $X=47300 $Y=-46365 $D=0
M124 238 67 GND GND NM L=1.8e-07 W=4.4e-07 $X=47300 $Y=9135 $D=0
M125 GND 264 69 GND NM L=1.8e-07 W=4.4e-07 $X=47600 $Y=-42665 $D=0
M126 GND 265 70 GND NM L=1.8e-07 W=4.4e-07 $X=47600 $Y=5435 $D=0
M127 GND 228 240 GND NM L=1.8e-07 W=4.4e-07 $X=47820 $Y=-29715 $D=0
M128 GND 229 241 GND NM L=1.8e-07 W=4.4e-07 $X=47820 $Y=-7515 $D=0
M129 GND 220 57 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-61710 $D=0
M130 GND 221 106 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-59910 $D=0
M131 GND 222 119 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-55090 $D=0
M132 GND 223 132 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-53290 $D=0
M133 GND 224 133 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=16280 $D=0
M134 GND 225 120 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=18080 $D=0
M135 GND 226 107 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=22900 $D=0
M136 GND 227 58 GND NM L=1.8e-07 W=2.2e-07 $X=47910 $Y=24700 $D=0
M137 245 200 GND GND NM L=1.8e-07 W=2.2e-07 $X=47940 $Y=-20365 $D=0
M138 242 59 GND GND NM L=1.8e-07 W=4.4e-07 $X=47940 $Y=-16765 $D=0
M139 GND 64 237 GND NM L=1.8e-07 W=4.4e-07 $X=48020 $Y=-46365 $D=0
M140 GND 230 233 GND NM L=1.8e-07 W=4.4e-07 $X=48020 $Y=-33415 $D=0
M141 GND 231 235 GND NM L=1.8e-07 W=4.4e-07 $X=48020 $Y=-3815 $D=0
M142 GND 65 238 GND NM L=1.8e-07 W=4.4e-07 $X=48020 $Y=9135 $D=0
M143 228 69 GND GND NM L=1.8e-07 W=2.2e-07 $X=48580 $Y=-29595 $D=0
M144 229 70 GND GND NM L=1.8e-07 W=2.2e-07 $X=48580 $Y=-7415 $D=0
M145 72 243 GND GND NM L=1.8e-07 W=4.4e-07 $X=48740 $Y=-46365 $D=0
M146 463 62 GND GND NM L=1.8e-07 W=4.4e-07 $X=48740 $Y=-33415 $D=0
M147 464 63 GND GND NM L=1.8e-07 W=4.4e-07 $X=48740 $Y=-3815 $D=0
M148 73 244 GND GND NM L=1.8e-07 W=4.4e-07 $X=48740 $Y=9135 $D=0
M149 230 69 463 GND NM L=1.8e-07 W=4.4e-07 $X=49170 $Y=-33415 $D=0
M150 231 70 464 GND NM L=1.8e-07 W=4.4e-07 $X=49170 $Y=-3815 $D=0
M151 GND 75 248 GND NM L=1.8e-07 W=4.4e-07 $X=49540 $Y=-42665 $D=0
M152 GND 76 251 GND NM L=1.8e-07 W=4.4e-07 $X=49540 $Y=5435 $D=0
M153 246 245 GND GND NM L=1.8e-07 W=4.4e-07 $X=49920 $Y=-20465 $D=0
M154 247 232 GND GND NM L=1.8e-07 W=4.4e-07 $X=49920 $Y=-16765 $D=0
M155 465 75 GND GND NM L=1.8e-07 W=4.4e-07 $X=50260 $Y=-42665 $D=0
M156 466 76 GND GND NM L=1.8e-07 W=4.4e-07 $X=50260 $Y=5435 $D=0
M157 Q6I 71 246 GND NM L=1.8e-07 W=4.4e-07 $X=50680 $Y=-20465 $D=0
M158 264 79 465 GND NM L=1.8e-07 W=4.4e-07 $X=50690 $Y=-42665 $D=0
M159 265 80 466 GND NM L=1.8e-07 W=4.4e-07 $X=50690 $Y=5435 $D=0
M160 GND 256 79 GND NM L=1.8e-07 W=2.2e-07 $X=50720 $Y=-46265 $D=0
M161 GND 257 80 GND NM L=1.8e-07 W=2.2e-07 $X=50720 $Y=9255 $D=0
M162 258 230 252 GND NM L=1.8e-07 W=4.4e-07 $X=51110 $Y=-33415 $D=0
M163 259 231 253 GND NM L=1.8e-07 W=4.4e-07 $X=51110 $Y=-3815 $D=0
M164 467 69 260 GND NM L=1.8e-07 W=4.4e-07 $X=51360 $Y=-29715 $D=0
M165 468 70 261 GND NM L=1.8e-07 W=4.4e-07 $X=51360 $Y=-7515 $D=0
M166 248 72 264 GND NM L=1.8e-07 W=4.4e-07 $X=51410 $Y=-42665 $D=0
M167 251 73 265 GND NM L=1.8e-07 W=4.4e-07 $X=51410 $Y=5435 $D=0
M168 GND 62 467 GND NM L=1.8e-07 W=4.4e-07 $X=51790 $Y=-29715 $D=0
M169 GND 63 468 GND NM L=1.8e-07 W=4.4e-07 $X=51790 $Y=-7515 $D=0
M170 GND 62 258 GND NM L=1.8e-07 W=4.4e-07 $X=51830 $Y=-33415 $D=0
M171 GND 63 259 GND NM L=1.8e-07 W=4.4e-07 $X=51830 $Y=-3815 $D=0
M172 GND 79 248 GND NM L=1.8e-07 W=4.4e-07 $X=52130 $Y=-42665 $D=0
M173 GND 80 251 GND NM L=1.8e-07 W=4.4e-07 $X=52130 $Y=5435 $D=0
M174 258 69 GND GND NM L=1.8e-07 W=4.4e-07 $X=52550 $Y=-33415 $D=0
M175 260 228 GND GND NM L=1.8e-07 W=2.2e-07 $X=52550 $Y=-29595 $D=0
M176 261 229 GND GND NM L=1.8e-07 W=2.2e-07 $X=52550 $Y=-7415 $D=0
M177 259 70 GND GND NM L=1.8e-07 W=4.4e-07 $X=52550 $Y=-3815 $D=0
M178 469 79 GND GND NM L=1.8e-07 W=4.4e-07 $X=52850 $Y=-42665 $D=0
M179 470 80 GND GND NM L=1.8e-07 W=4.4e-07 $X=52850 $Y=5435 $D=0
M180 471 75 469 GND NM L=1.8e-07 W=4.4e-07 $X=53280 $Y=-42665 $D=0
M181 472 76 470 GND NM L=1.8e-07 W=4.4e-07 $X=53280 $Y=5435 $D=0
M182 280 72 471 GND NM L=1.8e-07 W=4.4e-07 $X=53710 $Y=-42665 $D=0
M183 281 73 472 GND NM L=1.8e-07 W=4.4e-07 $X=53710 $Y=5435 $D=0
M184 276 264 280 GND NM L=1.8e-07 W=4.4e-07 $X=54430 $Y=-42665 $D=0
M185 279 265 281 GND NM L=1.8e-07 W=4.4e-07 $X=54430 $Y=5435 $D=0
M186 270 252 GND GND NM L=1.8e-07 W=4.4e-07 $X=54530 $Y=-33415 $D=0
M187 268 260 GND GND NM L=1.8e-07 W=4.4e-07 $X=54530 $Y=-29715 $D=0
M188 269 261 GND GND NM L=1.8e-07 W=4.4e-07 $X=54530 $Y=-7515 $D=0
M189 271 253 GND GND NM L=1.8e-07 W=4.4e-07 $X=54530 $Y=-3815 $D=0
M190 273 93 71 GND NM L=1.8e-07 W=4.4e-07 $X=54560 $Y=-20465 $D=0
M191 GND 60 274 GND NM L=1.8e-07 W=4.4e-07 $X=54570 $Y=-46365 $D=0
M192 GND 61 275 GND NM L=1.8e-07 W=4.4e-07 $X=54570 $Y=9135 $D=0
M193 GND 72 276 GND NM L=1.8e-07 W=4.4e-07 $X=55150 $Y=-42665 $D=0
M194 GND 73 279 GND NM L=1.8e-07 W=4.4e-07 $X=55150 $Y=5435 $D=0
M195 GND 262 273 GND NM L=1.8e-07 W=4.4e-07 $X=55280 $Y=-20465 $D=0
M196 84 81 268 GND NM L=1.8e-07 W=4.4e-07 $X=55290 $Y=-29715 $D=0
M197 74 82 269 GND NM L=1.8e-07 W=4.4e-07 $X=55290 $Y=-7515 $D=0
M198 GND 263 272 GND NM L=1.8e-07 W=4.4e-07 $X=55480 $Y=-16765 $D=0
M199 276 75 GND GND NM L=1.8e-07 W=4.4e-07 $X=55870 $Y=-42665 $D=0
M200 279 76 GND GND NM L=1.8e-07 W=4.4e-07 $X=55870 $Y=5435 $D=0
M201 262 84 GND GND NM L=1.8e-07 W=2.2e-07 $X=56040 $Y=-20365 $D=0
M202 473 74 GND GND NM L=1.8e-07 W=4.4e-07 $X=56200 $Y=-16765 $D=0
M203 GND 79 276 GND NM L=1.8e-07 W=4.4e-07 $X=56590 $Y=-42665 $D=0
M204 GND 80 279 GND NM L=1.8e-07 W=4.4e-07 $X=56590 $Y=5435 $D=0
M205 263 84 473 GND NM L=1.8e-07 W=4.4e-07 $X=56630 $Y=-16765 $D=0
M206 98 266 GND GND NM L=1.8e-07 W=2.2e-07 $X=57270 $Y=-46265 $D=0
M207 99 267 GND GND NM L=1.8e-07 W=2.2e-07 $X=57270 $Y=9255 $D=0
M208 86 280 GND GND NM L=1.8e-07 W=4.4e-07 $X=57310 $Y=-42665 $D=0
M209 87 281 GND GND NM L=1.8e-07 W=4.4e-07 $X=57310 $Y=5435 $D=0
M210 296 263 290 GND NM L=1.8e-07 W=4.4e-07 $X=58570 $Y=-16765 $D=0
M211 474 84 297 GND NM L=1.8e-07 W=4.4e-07 $X=58820 $Y=-20465 $D=0
M212 294 288 81 GND NM L=1.8e-07 W=4.4e-07 $X=59170 $Y=-29715 $D=0
M213 295 289 82 GND NM L=1.8e-07 W=4.4e-07 $X=59170 $Y=-7515 $D=0
M214 GND 320 88 GND NM L=1.8e-07 W=4.4e-07 $X=59250 $Y=-42665 $D=0
M215 GND 74 474 GND NM L=1.8e-07 W=4.4e-07 $X=59250 $Y=-20465 $D=0
M216 GND 321 89 GND NM L=1.8e-07 W=4.4e-07 $X=59250 $Y=5435 $D=0
M217 GND 298 75 GND NM L=1.8e-07 W=2.2e-07 $X=59290 $Y=-46265 $D=0
M218 GND 74 296 GND NM L=1.8e-07 W=4.4e-07 $X=59290 $Y=-16765 $D=0
M219 GND 299 76 GND NM L=1.8e-07 W=2.2e-07 $X=59290 $Y=9255 $D=0
M220 GND 282 294 GND NM L=1.8e-07 W=4.4e-07 $X=59890 $Y=-29715 $D=0
M221 GND 283 295 GND NM L=1.8e-07 W=4.4e-07 $X=59890 $Y=-7515 $D=0
M222 297 262 GND GND NM L=1.8e-07 W=2.2e-07 $X=60010 $Y=-20365 $D=0
M223 296 84 GND GND NM L=1.8e-07 W=4.4e-07 $X=60010 $Y=-16765 $D=0
M224 GND 284 291 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=-33415 $D=0
M225 GND 285 293 GND NM L=1.8e-07 W=4.4e-07 $X=60090 $Y=-3815 $D=0
M226 282 88 GND GND NM L=1.8e-07 W=2.2e-07 $X=60650 $Y=-29595 $D=0
M227 283 89 GND GND NM L=1.8e-07 W=2.2e-07 $X=60650 $Y=-7415 $D=0
M228 475 86 GND GND NM L=1.8e-07 W=4.4e-07 $X=60810 $Y=-33415 $D=0
M229 476 87 GND GND NM L=1.8e-07 W=4.4e-07 $X=60810 $Y=-3815 $D=0
M230 GND 96 304 GND NM L=1.8e-07 W=4.4e-07 $X=61190 $Y=-42665 $D=0
M231 GND 97 307 GND NM L=1.8e-07 W=4.4e-07 $X=61190 $Y=5435 $D=0
M232 284 88 475 GND NM L=1.8e-07 W=4.4e-07 $X=61240 $Y=-33415 $D=0
M233 285 89 476 GND NM L=1.8e-07 W=4.4e-07 $X=61240 $Y=-3815 $D=0
M234 477 96 GND GND NM L=1.8e-07 W=4.4e-07 $X=61910 $Y=-42665 $D=0
M235 478 97 GND GND NM L=1.8e-07 W=4.4e-07 $X=61910 $Y=5435 $D=0
M236 300 297 GND GND NM L=1.8e-07 W=4.4e-07 $X=61990 $Y=-20465 $D=0
M237 301 290 GND GND NM L=1.8e-07 W=4.4e-07 $X=61990 $Y=-16765 $D=0
M238 320 98 477 GND NM L=1.8e-07 W=4.4e-07 $X=62340 $Y=-42665 $D=0
M239 321 99 478 GND NM L=1.8e-07 W=4.4e-07 $X=62340 $Y=5435 $D=0
M240 Q5I 93 300 GND NM L=1.8e-07 W=4.4e-07 $X=62750 $Y=-20465 $D=0
M241 304 94 320 GND NM L=1.8e-07 W=4.4e-07 $X=63060 $Y=-42665 $D=0
M242 307 95 321 GND NM L=1.8e-07 W=4.4e-07 $X=63060 $Y=5435 $D=0
M243 GND 83 310 GND NM L=1.8e-07 W=4.4e-07 $X=63140 $Y=-46365 $D=0
M244 GND 85 311 GND NM L=1.8e-07 W=4.4e-07 $X=63140 $Y=9135 $D=0
M245 314 284 308 GND NM L=1.8e-07 W=4.4e-07 $X=63180 $Y=-33415 $D=0
M246 315 285 309 GND NM L=1.8e-07 W=4.4e-07 $X=63180 $Y=-3815 $D=0
M247 479 88 316 GND NM L=1.8e-07 W=4.4e-07 $X=63430 $Y=-29715 $D=0
M248 480 89 317 GND NM L=1.8e-07 W=4.4e-07 $X=63430 $Y=-7515 $D=0
M249 GND 98 304 GND NM L=1.8e-07 W=4.4e-07 $X=63780 $Y=-42665 $D=0
M250 GND 99 307 GND NM L=1.8e-07 W=4.4e-07 $X=63780 $Y=5435 $D=0
M251 GND 86 479 GND NM L=1.8e-07 W=4.4e-07 $X=63860 $Y=-29715 $D=0
M252 GND 87 480 GND NM L=1.8e-07 W=4.4e-07 $X=63860 $Y=-7515 $D=0
M253 GND 86 314 GND NM L=1.8e-07 W=4.4e-07 $X=63900 $Y=-33415 $D=0
M254 GND 87 315 GND NM L=1.8e-07 W=4.4e-07 $X=63900 $Y=-3815 $D=0
M255 481 98 GND GND NM L=1.8e-07 W=4.4e-07 $X=64500 $Y=-42665 $D=0
M256 482 99 GND GND NM L=1.8e-07 W=4.4e-07 $X=64500 $Y=5435 $D=0
M257 314 88 GND GND NM L=1.8e-07 W=4.4e-07 $X=64620 $Y=-33415 $D=0
M258 316 282 GND GND NM L=1.8e-07 W=2.2e-07 $X=64620 $Y=-29595 $D=0
M259 317 283 GND GND NM L=1.8e-07 W=2.2e-07 $X=64620 $Y=-7415 $D=0
M260 315 89 GND GND NM L=1.8e-07 W=4.4e-07 $X=64620 $Y=-3815 $D=0
M261 483 96 481 GND NM L=1.8e-07 W=4.4e-07 $X=64930 $Y=-42665 $D=0
M262 484 97 482 GND NM L=1.8e-07 W=4.4e-07 $X=64930 $Y=5435 $D=0
M263 332 94 483 GND NM L=1.8e-07 W=4.4e-07 $X=65360 $Y=-42665 $D=0
M264 333 95 484 GND NM L=1.8e-07 W=4.4e-07 $X=65360 $Y=5435 $D=0
M265 96 302 GND GND NM L=1.8e-07 W=2.2e-07 $X=65840 $Y=-46265 $D=0
M266 97 303 GND GND NM L=1.8e-07 W=2.2e-07 $X=65840 $Y=9255 $D=0
M267 328 320 332 GND NM L=1.8e-07 W=4.4e-07 $X=66080 $Y=-42665 $D=0
M268 331 321 333 GND NM L=1.8e-07 W=4.4e-07 $X=66080 $Y=5435 $D=0
M269 324 308 GND GND NM L=1.8e-07 W=4.4e-07 $X=66600 $Y=-33415 $D=0
M270 322 316 GND GND NM L=1.8e-07 W=4.4e-07 $X=66600 $Y=-29715 $D=0
M271 323 317 GND GND NM L=1.8e-07 W=4.4e-07 $X=66600 $Y=-7515 $D=0
M272 325 309 GND GND NM L=1.8e-07 W=4.4e-07 $X=66600 $Y=-3815 $D=0
M273 327 113 93 GND NM L=1.8e-07 W=4.4e-07 $X=66630 $Y=-20465 $D=0
M274 GND 94 328 GND NM L=1.8e-07 W=4.4e-07 $X=66800 $Y=-42665 $D=0
M275 GND 95 331 GND NM L=1.8e-07 W=4.4e-07 $X=66800 $Y=5435 $D=0
M276 GND 318 327 GND NM L=1.8e-07 W=4.4e-07 $X=67350 $Y=-20465 $D=0
M277 103 288 322 GND NM L=1.8e-07 W=4.4e-07 $X=67360 $Y=-29715 $D=0
M278 100 289 323 GND NM L=1.8e-07 W=4.4e-07 $X=67360 $Y=-7515 $D=0
M279 328 96 GND GND NM L=1.8e-07 W=4.4e-07 $X=67520 $Y=-42665 $D=0
M280 331 97 GND GND NM L=1.8e-07 W=4.4e-07 $X=67520 $Y=5435 $D=0
M281 GND 319 326 GND NM L=1.8e-07 W=4.4e-07 $X=67550 $Y=-16765 $D=0
M282 GND 356 94 GND NM L=1.8e-07 W=4.4e-07 $X=67820 $Y=-46365 $D=0
M283 GND 357 95 GND NM L=1.8e-07 W=4.4e-07 $X=67820 $Y=9135 $D=0
M284 318 103 GND GND NM L=1.8e-07 W=2.2e-07 $X=68110 $Y=-20365 $D=0
M285 GND 98 328 GND NM L=1.8e-07 W=4.4e-07 $X=68240 $Y=-42665 $D=0
M286 GND 99 331 GND NM L=1.8e-07 W=4.4e-07 $X=68240 $Y=5435 $D=0
M287 485 100 GND GND NM L=1.8e-07 W=4.4e-07 $X=68270 $Y=-16765 $D=0
M288 319 103 485 GND NM L=1.8e-07 W=4.4e-07 $X=68700 $Y=-16765 $D=0
M289 104 332 GND GND NM L=1.8e-07 W=4.4e-07 $X=68960 $Y=-42665 $D=0
M290 105 333 GND GND NM L=1.8e-07 W=4.4e-07 $X=68960 $Y=5435 $D=0
M291 GND 286 288 GND NM L=1.8e-07 W=2.2e-07 $X=69340 $Y=-33315 $D=0
M292 342 Q3I GND GND NM L=1.8e-07 W=2.2e-07 $X=69340 $Y=-29595 $D=0
M293 343 Q8I GND GND NM L=1.8e-07 W=2.2e-07 $X=69340 $Y=-7415 $D=0
M294 GND 287 289 GND NM L=1.8e-07 W=2.2e-07 $X=69340 $Y=-3695 $D=0
M295 GND 108 339 GND NM L=1.8e-07 W=4.4e-07 $X=69760 $Y=-46365 $D=0
M296 GND 109 340 GND NM L=1.8e-07 W=4.4e-07 $X=69760 $Y=9135 $D=0
M297 486 108 GND GND NM L=1.8e-07 W=4.4e-07 $X=70480 $Y=-46365 $D=0
M298 487 109 GND GND NM L=1.8e-07 W=4.4e-07 $X=70480 $Y=9135 $D=0
M299 344 319 336 GND NM L=1.8e-07 W=4.4e-07 $X=70640 $Y=-16765 $D=0
M300 488 103 345 GND NM L=1.8e-07 W=4.4e-07 $X=70890 $Y=-20465 $D=0
M301 356 38 486 GND NM L=1.8e-07 W=4.4e-07 $X=70910 $Y=-46365 $D=0
M302 357 39 487 GND NM L=1.8e-07 W=4.4e-07 $X=70910 $Y=9135 $D=0
M303 GND 346 101 GND NM L=1.8e-07 W=2.2e-07 $X=70940 $Y=-42545 $D=0
M304 GND 347 102 GND NM L=1.8e-07 W=2.2e-07 $X=70940 $Y=5535 $D=0
M305 334 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=71320 $Y=-29715 $D=0
M306 GND 100 488 GND NM L=1.8e-07 W=4.4e-07 $X=71320 $Y=-20465 $D=0
M307 335 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=71320 $Y=-7515 $D=0
M308 GND 100 344 GND NM L=1.8e-07 W=4.4e-07 $X=71360 $Y=-16765 $D=0
M309 339 106 356 GND NM L=1.8e-07 W=4.4e-07 $X=71630 $Y=-46365 $D=0
M310 340 107 357 GND NM L=1.8e-07 W=4.4e-07 $X=71630 $Y=9135 $D=0
M311 GND 342 334 GND NM L=1.8e-07 W=4.4e-07 $X=72040 $Y=-29715 $D=0
M312 GND 343 335 GND NM L=1.8e-07 W=4.4e-07 $X=72040 $Y=-7515 $D=0
M313 345 318 GND GND NM L=1.8e-07 W=2.2e-07 $X=72080 $Y=-20365 $D=0
M314 344 103 GND GND NM L=1.8e-07 W=4.4e-07 $X=72080 $Y=-16765 $D=0
M315 GND 38 339 GND NM L=1.8e-07 W=4.4e-07 $X=72350 $Y=-46365 $D=0
M316 GND 39 340 GND NM L=1.8e-07 W=4.4e-07 $X=72350 $Y=9135 $D=0
M317 489 334 GND GND NM L=1.8e-07 W=4.4e-07 $X=72760 $Y=-29715 $D=0
M318 490 335 GND GND NM L=1.8e-07 W=4.4e-07 $X=72760 $Y=-7515 $D=0
M319 491 38 GND GND NM L=1.8e-07 W=4.4e-07 $X=73070 $Y=-46365 $D=0
M320 492 39 GND GND NM L=1.8e-07 W=4.4e-07 $X=73070 $Y=9135 $D=0
M321 GND 101 352 GND NM L=1.8e-07 W=4.4e-07 $X=73190 $Y=-33415 $D=0
M322 350 CLK 489 GND NM L=1.8e-07 W=4.4e-07 $X=73190 $Y=-29715 $D=0
M323 351 CLK 490 GND NM L=1.8e-07 W=4.4e-07 $X=73190 $Y=-7515 $D=0
M324 GND 102 353 GND NM L=1.8e-07 W=4.4e-07 $X=73190 $Y=-3815 $D=0
M325 493 108 491 GND NM L=1.8e-07 W=4.4e-07 $X=73500 $Y=-46365 $D=0
M326 494 109 492 GND NM L=1.8e-07 W=4.4e-07 $X=73500 $Y=9135 $D=0
M327 370 106 493 GND NM L=1.8e-07 W=4.4e-07 $X=73930 $Y=-46365 $D=0
M328 371 107 494 GND NM L=1.8e-07 W=4.4e-07 $X=73930 $Y=9135 $D=0
M329 354 345 GND GND NM L=1.8e-07 W=4.4e-07 $X=74060 $Y=-20465 $D=0
M330 355 336 GND GND NM L=1.8e-07 W=4.4e-07 $X=74060 $Y=-16765 $D=0
M331 365 356 370 GND NM L=1.8e-07 W=4.4e-07 $X=74650 $Y=-46365 $D=0
M332 366 357 371 GND NM L=1.8e-07 W=4.4e-07 $X=74650 $Y=9135 $D=0
M333 GND 114 362 GND NM L=1.8e-07 W=4.4e-07 $X=74790 $Y=-42665 $D=0
M334 GND 115 363 GND NM L=1.8e-07 W=4.4e-07 $X=74790 $Y=5435 $D=0
M335 Q4I 113 354 GND NM L=1.8e-07 W=4.4e-07 $X=74820 $Y=-20465 $D=0
M336 495 CLK Q3 GND NM L=1.8e-07 W=4.4e-07 $X=75130 $Y=-29715 $D=0
M337 496 CLK Q8 GND NM L=1.8e-07 W=4.4e-07 $X=75130 $Y=-7515 $D=0
M338 GND 106 365 GND NM L=1.8e-07 W=4.4e-07 $X=75370 $Y=-46365 $D=0
M339 GND 107 366 GND NM L=1.8e-07 W=4.4e-07 $X=75370 $Y=9135 $D=0
M340 GND 350 495 GND NM L=1.8e-07 W=4.4e-07 $X=75560 $Y=-29715 $D=0
M341 GND 351 496 GND NM L=1.8e-07 W=4.4e-07 $X=75560 $Y=-7515 $D=0
M342 121 348 GND GND NM L=1.8e-07 W=2.2e-07 $X=75890 $Y=-33315 $D=0
M343 118 349 GND GND NM L=1.8e-07 W=2.2e-07 $X=75890 $Y=-3695 $D=0
M344 365 108 GND GND NM L=1.8e-07 W=4.4e-07 $X=76090 $Y=-46365 $D=0
M345 366 109 GND GND NM L=1.8e-07 W=4.4e-07 $X=76090 $Y=9135 $D=0
M346 INVQ3 Q3 GND GND NM L=1.8e-07 W=4.4e-07 $X=76280 $Y=-29715 $D=0
M347 INVQ8 Q8 GND GND NM L=1.8e-07 W=4.4e-07 $X=76280 $Y=-7515 $D=0
M348 GND 38 365 GND NM L=1.8e-07 W=4.4e-07 $X=76810 $Y=-46365 $D=0
M349 GND 39 366 GND NM L=1.8e-07 W=4.4e-07 $X=76810 $Y=9135 $D=0
M350 125 358 GND GND NM L=1.8e-07 W=2.2e-07 $X=77490 $Y=-42545 $D=0
M351 124 359 GND GND NM L=1.8e-07 W=2.2e-07 $X=77490 $Y=5535 $D=0
M352 111 370 GND GND NM L=1.8e-07 W=4.4e-07 $X=77530 $Y=-46365 $D=0
M353 112 371 GND GND NM L=1.8e-07 W=4.4e-07 $X=77530 $Y=9135 $D=0
M354 378 Q2I GND GND NM L=1.8e-07 W=2.2e-07 $X=78260 $Y=-29595 $D=0
M355 379 Q7I GND GND NM L=1.8e-07 W=2.2e-07 $X=78260 $Y=-7415 $D=0
M356 375 123 113 GND NM L=1.8e-07 W=4.4e-07 $X=78700 $Y=-20465 $D=0
M357 GND 372 375 GND NM L=1.8e-07 W=4.4e-07 $X=79420 $Y=-20465 $D=0
M358 GND 380 114 GND NM L=1.8e-07 W=2.2e-07 $X=79510 $Y=-46265 $D=0
M359 GND 381 115 GND NM L=1.8e-07 W=2.2e-07 $X=79510 $Y=9255 $D=0
M360 GND 373 374 GND NM L=1.8e-07 W=4.4e-07 $X=79620 $Y=-16765 $D=0
M361 372 121 GND GND NM L=1.8e-07 W=2.2e-07 $X=80180 $Y=-20365 $D=0
M362 376 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=80240 $Y=-29715 $D=0
M363 377 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=80240 $Y=-7515 $D=0
M364 497 118 GND GND NM L=1.8e-07 W=4.4e-07 $X=80340 $Y=-16765 $D=0
M365 373 121 497 GND NM L=1.8e-07 W=4.4e-07 $X=80770 $Y=-16765 $D=0
M366 GND 378 376 GND NM L=1.8e-07 W=4.4e-07 $X=80960 $Y=-29715 $D=0
M367 GND 379 377 GND NM L=1.8e-07 W=4.4e-07 $X=80960 $Y=-7515 $D=0
M368 498 376 GND GND NM L=1.8e-07 W=4.4e-07 $X=81680 $Y=-29715 $D=0
M369 499 377 GND GND NM L=1.8e-07 W=4.4e-07 $X=81680 $Y=-7515 $D=0
M370 382 CLK 498 GND NM L=1.8e-07 W=4.4e-07 $X=82110 $Y=-29715 $D=0
M371 383 CLK 499 GND NM L=1.8e-07 W=4.4e-07 $X=82110 $Y=-7515 $D=0
M372 392 373 386 GND NM L=1.8e-07 W=4.4e-07 $X=82710 $Y=-16765 $D=0
M373 500 121 393 GND NM L=1.8e-07 W=4.4e-07 $X=82960 $Y=-20465 $D=0
M374 GND 116 390 GND NM L=1.8e-07 W=4.4e-07 $X=83360 $Y=-46365 $D=0
M375 GND 117 391 GND NM L=1.8e-07 W=4.4e-07 $X=83360 $Y=9135 $D=0
M376 GND 118 500 GND NM L=1.8e-07 W=4.4e-07 $X=83390 $Y=-20465 $D=0
M377 GND 118 392 GND NM L=1.8e-07 W=4.4e-07 $X=83430 $Y=-16765 $D=0
M378 501 CLK Q2 GND NM L=1.8e-07 W=4.4e-07 $X=84050 $Y=-29715 $D=0
M379 502 CLK Q7 GND NM L=1.8e-07 W=4.4e-07 $X=84050 $Y=-7515 $D=0
M380 393 372 GND GND NM L=1.8e-07 W=2.2e-07 $X=84150 $Y=-20365 $D=0
M381 392 121 GND GND NM L=1.8e-07 W=4.4e-07 $X=84150 $Y=-16765 $D=0
M382 GND 382 501 GND NM L=1.8e-07 W=4.4e-07 $X=84480 $Y=-29715 $D=0
M383 GND 383 502 GND NM L=1.8e-07 W=4.4e-07 $X=84480 $Y=-7515 $D=0
M384 INVQ2 Q2 GND GND NM L=1.8e-07 W=4.4e-07 $X=85200 $Y=-29715 $D=0
M385 INVQ7 Q7 GND GND NM L=1.8e-07 W=4.4e-07 $X=85200 $Y=-7515 $D=0
M386 131 384 GND GND NM L=1.8e-07 W=2.2e-07 $X=86060 $Y=-46265 $D=0
M387 128 385 GND GND NM L=1.8e-07 W=2.2e-07 $X=86060 $Y=9255 $D=0
M388 396 393 GND GND NM L=1.8e-07 W=4.4e-07 $X=86130 $Y=-20465 $D=0
M389 397 386 GND GND NM L=1.8e-07 W=4.4e-07 $X=86130 $Y=-16765 $D=0
M390 Q3I 123 396 GND NM L=1.8e-07 W=4.4e-07 $X=86890 $Y=-20465 $D=0
M391 402 Q1I GND GND NM L=1.8e-07 W=2.2e-07 $X=87180 $Y=-29595 $D=0
M392 403 Q6I GND GND NM L=1.8e-07 W=2.2e-07 $X=87180 $Y=-7415 $D=0
M393 398 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=89160 $Y=-29715 $D=0
M394 399 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=89160 $Y=-7515 $D=0
M395 GND 402 398 GND NM L=1.8e-07 W=4.4e-07 $X=89880 $Y=-29715 $D=0
M396 GND 403 399 GND NM L=1.8e-07 W=4.4e-07 $X=89880 $Y=-7515 $D=0
M397 503 398 GND GND NM L=1.8e-07 W=4.4e-07 $X=90600 $Y=-29715 $D=0
M398 504 399 GND GND NM L=1.8e-07 W=4.4e-07 $X=90600 $Y=-7515 $D=0
M399 405 127 123 GND NM L=1.8e-07 W=4.4e-07 $X=90770 $Y=-20465 $D=0
M400 406 CLK 503 GND NM L=1.8e-07 W=4.4e-07 $X=91030 $Y=-29715 $D=0
M401 407 CLK 504 GND NM L=1.8e-07 W=4.4e-07 $X=91030 $Y=-7515 $D=0
M402 GND 400 405 GND NM L=1.8e-07 W=4.4e-07 $X=91490 $Y=-20465 $D=0
M403 GND 401 404 GND NM L=1.8e-07 W=4.4e-07 $X=91690 $Y=-16765 $D=0
M404 400 125 GND GND NM L=1.8e-07 W=2.2e-07 $X=92250 $Y=-20365 $D=0
M405 505 124 GND GND NM L=1.8e-07 W=4.4e-07 $X=92410 $Y=-16765 $D=0
M406 401 125 505 GND NM L=1.8e-07 W=4.4e-07 $X=92840 $Y=-16765 $D=0
M407 506 CLK Q1 GND NM L=1.8e-07 W=4.4e-07 $X=92970 $Y=-29715 $D=0
M408 507 CLK Q6 GND NM L=1.8e-07 W=4.4e-07 $X=92970 $Y=-7515 $D=0
M409 GND 406 506 GND NM L=1.8e-07 W=4.4e-07 $X=93400 $Y=-29715 $D=0
M410 GND 407 507 GND NM L=1.8e-07 W=4.4e-07 $X=93400 $Y=-7515 $D=0
M411 INVQ1 Q1 GND GND NM L=1.8e-07 W=4.4e-07 $X=94120 $Y=-29715 $D=0
M412 INVQ6 Q6 GND GND NM L=1.8e-07 W=4.4e-07 $X=94120 $Y=-7515 $D=0
M413 414 401 412 GND NM L=1.8e-07 W=4.4e-07 $X=94780 $Y=-16765 $D=0
M414 508 125 415 GND NM L=1.8e-07 W=4.4e-07 $X=95030 $Y=-20465 $D=0
M415 GND 124 508 GND NM L=1.8e-07 W=4.4e-07 $X=95460 $Y=-20465 $D=0
M416 GND 124 414 GND NM L=1.8e-07 W=4.4e-07 $X=95500 $Y=-16765 $D=0
M417 420 Q0I GND GND NM L=1.8e-07 W=2.2e-07 $X=96100 $Y=-29595 $D=0
M418 421 Q5I GND GND NM L=1.8e-07 W=2.2e-07 $X=96100 $Y=-7415 $D=0
M419 415 400 GND GND NM L=1.8e-07 W=2.2e-07 $X=96220 $Y=-20365 $D=0
M420 414 125 GND GND NM L=1.8e-07 W=4.4e-07 $X=96220 $Y=-16765 $D=0
M421 416 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=98080 $Y=-29715 $D=0
M422 417 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=98080 $Y=-7515 $D=0
M423 418 415 GND GND NM L=1.8e-07 W=4.4e-07 $X=98200 $Y=-20465 $D=0
M424 419 412 GND GND NM L=1.8e-07 W=4.4e-07 $X=98200 $Y=-16765 $D=0
M425 GND 420 416 GND NM L=1.8e-07 W=4.4e-07 $X=98800 $Y=-29715 $D=0
M426 GND 421 417 GND NM L=1.8e-07 W=4.4e-07 $X=98800 $Y=-7515 $D=0
M427 Q2I 127 418 GND NM L=1.8e-07 W=4.4e-07 $X=98960 $Y=-20465 $D=0
M428 509 416 GND GND NM L=1.8e-07 W=4.4e-07 $X=99520 $Y=-29715 $D=0
M429 510 417 GND GND NM L=1.8e-07 W=4.4e-07 $X=99520 $Y=-7515 $D=0
M430 422 CLK 509 GND NM L=1.8e-07 W=4.4e-07 $X=99950 $Y=-29715 $D=0
M431 423 CLK 510 GND NM L=1.8e-07 W=4.4e-07 $X=99950 $Y=-7515 $D=0
M432 511 CLK Q0 GND NM L=1.8e-07 W=4.4e-07 $X=101890 $Y=-29715 $D=0
M433 512 CLK Q5 GND NM L=1.8e-07 W=4.4e-07 $X=101890 $Y=-7515 $D=0
M434 GND 422 511 GND NM L=1.8e-07 W=4.4e-07 $X=102320 $Y=-29715 $D=0
M435 GND 423 512 GND NM L=1.8e-07 W=4.4e-07 $X=102320 $Y=-7515 $D=0
M436 433 429 127 GND NM L=1.8e-07 W=4.4e-07 $X=102840 $Y=-20465 $D=0
M437 INVQ0 Q0 GND GND NM L=1.8e-07 W=4.4e-07 $X=103040 $Y=-29715 $D=0
M438 INVQ5 Q5 GND GND NM L=1.8e-07 W=4.4e-07 $X=103040 $Y=-7515 $D=0
M439 GND 424 433 GND NM L=1.8e-07 W=4.4e-07 $X=103560 $Y=-20465 $D=0
M440 GND 425 430 GND NM L=1.8e-07 W=4.4e-07 $X=103760 $Y=-16765 $D=0
M441 424 131 GND GND NM L=1.8e-07 W=2.2e-07 $X=104320 $Y=-20365 $D=0
M442 513 128 GND GND NM L=1.8e-07 W=4.4e-07 $X=104480 $Y=-16765 $D=0
M443 425 131 513 GND NM L=1.8e-07 W=4.4e-07 $X=104910 $Y=-16765 $D=0
M444 436 Q4I GND GND NM L=1.8e-07 W=2.2e-07 $X=105020 $Y=-7415 $D=0
M445 438 425 435 GND NM L=1.8e-07 W=4.4e-07 $X=106850 $Y=-16765 $D=0
M446 434 RST GND GND NM L=1.8e-07 W=4.4e-07 $X=107000 $Y=-7515 $D=0
M447 514 131 439 GND NM L=1.8e-07 W=4.4e-07 $X=107100 $Y=-20465 $D=0
M448 GND 128 514 GND NM L=1.8e-07 W=4.4e-07 $X=107530 $Y=-20465 $D=0
M449 GND 128 438 GND NM L=1.8e-07 W=4.4e-07 $X=107570 $Y=-16765 $D=0
M450 GND 436 434 GND NM L=1.8e-07 W=4.4e-07 $X=107720 $Y=-7515 $D=0
M451 439 424 GND GND NM L=1.8e-07 W=2.2e-07 $X=108290 $Y=-20365 $D=0
M452 438 131 GND GND NM L=1.8e-07 W=4.4e-07 $X=108290 $Y=-16765 $D=0
M453 515 434 GND GND NM L=1.8e-07 W=4.4e-07 $X=108440 $Y=-7515 $D=0
M454 440 CLK 515 GND NM L=1.8e-07 W=4.4e-07 $X=108870 $Y=-7515 $D=0
M455 441 439 GND GND NM L=1.8e-07 W=4.4e-07 $X=110270 $Y=-20465 $D=0
M456 442 435 GND GND NM L=1.8e-07 W=4.4e-07 $X=110270 $Y=-16765 $D=0
M457 516 CLK Q4 GND NM L=1.8e-07 W=4.4e-07 $X=110810 $Y=-7515 $D=0
M458 Q1I 429 441 GND NM L=1.8e-07 W=4.4e-07 $X=111030 $Y=-20465 $D=0
M459 GND 440 516 GND NM L=1.8e-07 W=4.4e-07 $X=111240 $Y=-7515 $D=0
M460 INVQ4 Q4 GND GND NM L=1.8e-07 W=4.4e-07 $X=111960 $Y=-7515 $D=0
M461 GND 428 429 GND NM L=1.8e-07 W=2.2e-07 $X=113010 $Y=-16645 $D=0
M462 GND 132 446 GND NM L=1.8e-07 W=4.4e-07 $X=116860 $Y=-16765 $D=0
M463 Q0I 445 GND GND NM L=1.8e-07 W=2.2e-07 $X=119560 $Y=-16645 $D=0
M464 134 37 Q8I VDD PM L=1.8e-07 W=4.4e-07 $X=30540 $Y=-13320 $D=4
M465 144 16 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-49810 $D=4
M466 18 14 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-39220 $D=4
M467 18 21 27 VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-36860 $D=4
M468 19 22 20 VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=-370 $D=4
M469 19 15 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=1990 $D=4
M470 145 17 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=31260 $Y=12580 $D=4
M471 VDD 146 135 VDD PM L=1.8e-07 W=8.8e-07 $X=31340 $Y=-23910 $D=4
M472 147 20 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=32060 $Y=-13320 $D=4
M473 146 20 517 VDD PM L=1.8e-07 W=8.8e-07 $X=32490 $Y=-23910 $D=4
M474 83 139 A0 VDD PM L=1.8e-07 W=2.2e-07 $X=32560 $Y=-51950 $D=4
M475 85 140 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=32560 $Y=14940 $D=4
M476 VDD 27 147 VDD PM L=1.8e-07 W=4.4e-07 $X=32780 $Y=-13320 $D=4
M477 GND B3 25 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-63050 $D=4
M478 GND B3 16 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-58570 $D=4
M479 GND B3 66 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-56430 $D=4
M480 GND B3 83 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=-51950 $D=4
M481 GND X3 85 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=14940 $D=4
M482 GND X3 67 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=19420 $D=4
M483 GND X3 17 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=21560 $D=4
M484 GND X3 26 VDD PM L=1.8e-07 W=2.2e-07 $X=33360 $Y=26040 $D=4
M485 152 144 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=33920 $Y=-49810 $D=4
M486 153 18 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=33920 $Y=-39220 $D=4
M487 154 19 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=33920 $Y=1990 $D=4
M488 155 145 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=33920 $Y=12580 $D=4
M489 158 147 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=34720 $Y=-13320 $D=4
M490 VDD 25 518 VDD PM L=1.8e-07 W=8.8e-07 $X=35110 $Y=-39660 $D=4
M491 VDD 26 519 VDD PM L=1.8e-07 W=8.8e-07 $X=35110 $Y=1990 $D=4
M492 163 55 23 VDD PM L=1.8e-07 W=4.4e-07 $X=35150 $Y=-36860 $D=4
M493 164 20 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=35150 $Y=-23910 $D=4
M494 165 56 24 VDD PM L=1.8e-07 W=4.4e-07 $X=35150 $Y=-370 $D=4
M495 166 43 23 VDD PM L=1.8e-07 W=4.4e-07 $X=35190 $Y=-26270 $D=4
M496 171 B2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=35390 $Y=-52050 $D=4
M497 172 X2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=35390 $Y=14820 $D=4
M498 520 20 158 VDD PM L=1.8e-07 W=8.8e-07 $X=35480 $Y=-13760 $D=4
M499 177 146 164 VDD PM L=1.8e-07 W=8.8e-07 $X=35870 $Y=-23910 $D=4
M500 VDD 148 166 VDD PM L=1.8e-07 W=8.8e-07 $X=35950 $Y=-26710 $D=4
M501 VDD 149 167 VDD PM L=1.8e-07 W=8.8e-07 $X=35950 $Y=-10960 $D=4
M502 150 28 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=36670 $Y=-36860 $D=4
M503 521 33 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=36670 $Y=-10960 $D=4
M504 151 29 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=36670 $Y=-370 $D=4
M505 148 28 522 VDD PM L=1.8e-07 W=8.8e-07 $X=37100 $Y=-26710 $D=4
M506 VDD 32 150 VDD PM L=1.8e-07 W=4.4e-07 $X=37390 $Y=-36860 $D=4
M507 VDD 33 151 VDD PM L=1.8e-07 W=4.4e-07 $X=37390 $Y=-370 $D=4
M508 108 171 A0 VDD PM L=1.8e-07 W=2.2e-07 $X=37410 $Y=-51950 $D=4
M509 109 172 Y0 VDD PM L=1.8e-07 W=2.2e-07 $X=37410 $Y=14940 $D=4
M510 179 158 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=37850 $Y=-13760 $D=4
M511 GND B2 30 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-63050 $D=4
M512 GND B2 64 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-58570 $D=4
M513 GND B2 91 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-56430 $D=4
M514 GND B2 108 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=-51950 $D=4
M515 GND X2 109 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=14940 $D=4
M516 GND X2 92 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=19420 $D=4
M517 GND X2 65 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=21560 $D=4
M518 GND X2 31 VDD PM L=1.8e-07 W=2.2e-07 $X=38210 $Y=26040 $D=4
M519 Q7I 36 178 VDD PM L=1.8e-07 W=4.4e-07 $X=38570 $Y=-23910 $D=4
M520 Q7I 37 179 VDD PM L=1.8e-07 W=4.4e-07 $X=38610 $Y=-13320 $D=4
M521 VDD 218 34 VDD PM L=1.8e-07 W=8.8e-07 $X=39030 $Y=-49810 $D=4
M522 VDD 219 35 VDD PM L=1.8e-07 W=8.8e-07 $X=39030 $Y=12140 $D=4
M523 VDD 32 184 VDD PM L=1.8e-07 W=8.8e-07 $X=39040 $Y=-26710 $D=4
M524 182 150 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=39330 $Y=-36860 $D=4
M525 183 151 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=39330 $Y=-370 $D=4
M526 184 28 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=39760 $Y=-26710 $D=4
M527 185 29 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=39760 $Y=-10960 $D=4
M528 188 34 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=39830 $Y=-39220 $D=4
M529 189 35 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=39830 $Y=1990 $D=4
M530 VDD 32 523 VDD PM L=1.8e-07 W=8.8e-07 $X=40520 $Y=-36860 $D=4
M531 VDD 33 524 VDD PM L=1.8e-07 W=8.8e-07 $X=40520 $Y=-810 $D=4
M532 VDD 40 188 VDD PM L=1.8e-07 W=4.4e-07 $X=40550 $Y=-39220 $D=4
M533 VDD 41 189 VDD PM L=1.8e-07 W=4.4e-07 $X=40550 $Y=1990 $D=4
M534 201 71 36 VDD PM L=1.8e-07 W=4.4e-07 $X=40660 $Y=-13320 $D=4
M535 200 68 36 VDD PM L=1.8e-07 W=4.4e-07 $X=40710 $Y=-23910 $D=4
M536 VDD 66 210 VDD PM L=1.8e-07 W=8.8e-07 $X=40970 $Y=-49810 $D=4
M537 VDD 67 213 VDD PM L=1.8e-07 W=8.8e-07 $X=40970 $Y=12140 $D=4
M538 525 66 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41690 $Y=-49810 $D=4
M539 526 67 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=41690 $Y=12140 $D=4
M540 218 64 525 VDD PM L=1.8e-07 W=8.8e-07 $X=42120 $Y=-49810 $D=4
M541 219 65 526 VDD PM L=1.8e-07 W=8.8e-07 $X=42120 $Y=12140 $D=4
M542 202 198 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42420 $Y=-26710 $D=4
M543 203 199 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42420 $Y=-10960 $D=4
M544 204 182 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42460 $Y=-36860 $D=4
M545 205 183 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=42460 $Y=-810 $D=4
M546 208 188 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=42490 $Y=-39220 $D=4
M547 209 189 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=42490 $Y=1990 $D=4
M548 206 71 37 VDD PM L=1.8e-07 W=4.4e-07 $X=42610 $Y=-13320 $D=4
M549 210 53 218 VDD PM L=1.8e-07 W=8.8e-07 $X=42840 $Y=-49810 $D=4
M550 213 54 219 VDD PM L=1.8e-07 W=8.8e-07 $X=42840 $Y=12140 $D=4
M551 GND B1 53 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-63050 $D=4
M552 GND B1 60 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-58570 $D=4
M553 GND B1 38 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-56430 $D=4
M554 GND B1 116 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=-51950 $D=4
M555 GND X1 117 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=14940 $D=4
M556 GND X1 39 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=19420 $D=4
M557 GND X1 61 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=21560 $D=4
M558 GND X1 54 VDD PM L=1.8e-07 W=2.2e-07 $X=43060 $Y=26040 $D=4
M559 59 43 202 VDD PM L=1.8e-07 W=4.4e-07 $X=43180 $Y=-26270 $D=4
M560 42 44 203 VDD PM L=1.8e-07 W=4.4e-07 $X=43180 $Y=-10960 $D=4
M561 59 55 204 VDD PM L=1.8e-07 W=4.4e-07 $X=43220 $Y=-36860 $D=4
M562 42 56 205 VDD PM L=1.8e-07 W=4.4e-07 $X=43220 $Y=-370 $D=4
M563 VDD 200 207 VDD PM L=1.8e-07 W=8.8e-07 $X=43410 $Y=-23910 $D=4
M564 VDD 64 210 VDD PM L=1.8e-07 W=8.8e-07 $X=43560 $Y=-49810 $D=4
M565 VDD 65 213 VDD PM L=1.8e-07 W=8.8e-07 $X=43560 $Y=12140 $D=4
M566 VDD 40 527 VDD PM L=1.8e-07 W=8.8e-07 $X=43680 $Y=-39660 $D=4
M567 VDD 41 528 VDD PM L=1.8e-07 W=8.8e-07 $X=43680 $Y=1990 $D=4
M568 201 42 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=44130 $Y=-13320 $D=4
M569 529 64 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44280 $Y=-49810 $D=4
M570 530 65 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=44280 $Y=12140 $D=4
M571 531 66 529 VDD PM L=1.8e-07 W=8.8e-07 $X=44710 $Y=-49810 $D=4
M572 532 67 530 VDD PM L=1.8e-07 W=8.8e-07 $X=44710 $Y=12140 $D=4
M573 243 53 531 VDD PM L=1.8e-07 W=8.8e-07 $X=45140 $Y=-49810 $D=4
M574 244 54 532 VDD PM L=1.8e-07 W=8.8e-07 $X=45140 $Y=12140 $D=4
M575 230 81 43 VDD PM L=1.8e-07 W=4.4e-07 $X=45270 $Y=-36860 $D=4
M576 231 82 44 VDD PM L=1.8e-07 W=4.4e-07 $X=45270 $Y=-370 $D=4
M577 228 77 43 VDD PM L=1.8e-07 W=4.4e-07 $X=45320 $Y=-26270 $D=4
M578 229 78 44 VDD PM L=1.8e-07 W=4.4e-07 $X=45320 $Y=-10960 $D=4
M579 236 218 243 VDD PM L=1.8e-07 W=8.8e-07 $X=45860 $Y=-49810 $D=4
M580 239 219 244 VDD PM L=1.8e-07 W=8.8e-07 $X=45860 $Y=12140 $D=4
M581 VDD 53 236 VDD PM L=1.8e-07 W=8.8e-07 $X=46580 $Y=-49810 $D=4
M582 VDD 54 239 VDD PM L=1.8e-07 W=8.8e-07 $X=46580 $Y=12140 $D=4
M583 232 201 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=46790 $Y=-13320 $D=4
M584 233 81 55 VDD PM L=1.8e-07 W=4.4e-07 $X=47220 $Y=-36860 $D=4
M585 234 42 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=47220 $Y=-23910 $D=4
M586 235 82 56 VDD PM L=1.8e-07 W=4.4e-07 $X=47220 $Y=-370 $D=4
M587 240 77 55 VDD PM L=1.8e-07 W=4.4e-07 $X=47260 $Y=-26270 $D=4
M588 236 66 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=47300 $Y=-49810 $D=4
M589 239 67 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=47300 $Y=12140 $D=4
M590 533 42 232 VDD PM L=1.8e-07 W=8.8e-07 $X=47550 $Y=-13760 $D=4
M591 VDD 264 69 VDD PM L=1.8e-07 W=8.8e-07 $X=47600 $Y=-39660 $D=4
M592 VDD 265 70 VDD PM L=1.8e-07 W=8.8e-07 $X=47600 $Y=1990 $D=4
M593 GND B0 57 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-63050 $D=4
M594 GND B0 106 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-58570 $D=4
M595 GND B0 119 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-56430 $D=4
M596 GND B0 132 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=-51950 $D=4
M597 GND X0 133 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=14940 $D=4
M598 GND X0 120 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=19420 $D=4
M599 GND X0 107 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=21560 $D=4
M600 GND X0 58 VDD PM L=1.8e-07 W=2.2e-07 $X=47910 $Y=26040 $D=4
M601 VDD 59 533 VDD PM L=1.8e-07 W=8.8e-07 $X=47980 $Y=-13760 $D=4
M602 VDD 64 236 VDD PM L=1.8e-07 W=8.8e-07 $X=48020 $Y=-49810 $D=4
M603 VDD 228 240 VDD PM L=1.8e-07 W=8.8e-07 $X=48020 $Y=-26710 $D=4
M604 VDD 229 241 VDD PM L=1.8e-07 W=8.8e-07 $X=48020 $Y=-10960 $D=4
M605 VDD 65 239 VDD PM L=1.8e-07 W=8.8e-07 $X=48020 $Y=12140 $D=4
M606 72 243 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48740 $Y=-49810 $D=4
M607 230 62 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=48740 $Y=-36860 $D=4
M608 534 69 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48740 $Y=-26710 $D=4
M609 231 63 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=48740 $Y=-370 $D=4
M610 73 244 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=48740 $Y=12140 $D=4
M611 229 63 535 VDD PM L=1.8e-07 W=8.8e-07 $X=49170 $Y=-10960 $D=4
M612 VDD 75 249 VDD PM L=1.8e-07 W=8.8e-07 $X=49540 $Y=-39660 $D=4
M613 VDD 76 250 VDD PM L=1.8e-07 W=8.8e-07 $X=49540 $Y=1990 $D=4
M614 246 245 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=49880 $Y=-23910 $D=4
M615 536 75 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50260 $Y=-39660 $D=4
M616 537 76 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=50260 $Y=1990 $D=4
M617 Q6I 68 246 VDD PM L=1.8e-07 W=4.4e-07 $X=50640 $Y=-23910 $D=4
M618 Q6I 71 247 VDD PM L=1.8e-07 W=4.4e-07 $X=50680 $Y=-13320 $D=4
M619 264 79 536 VDD PM L=1.8e-07 W=8.8e-07 $X=50690 $Y=-39660 $D=4
M620 265 80 537 VDD PM L=1.8e-07 W=8.8e-07 $X=50690 $Y=1990 $D=4
M621 VDD 70 255 VDD PM L=1.8e-07 W=8.8e-07 $X=51110 $Y=-10960 $D=4
M622 252 230 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=51400 $Y=-36860 $D=4
M623 253 231 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=51400 $Y=-370 $D=4
M624 249 72 264 VDD PM L=1.8e-07 W=8.8e-07 $X=51410 $Y=-39660 $D=4
M625 250 73 265 VDD PM L=1.8e-07 W=8.8e-07 $X=51410 $Y=1990 $D=4
M626 256 60 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=51480 $Y=-49810 $D=4
M627 257 61 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=51480 $Y=12580 $D=4
M628 254 62 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=51830 $Y=-26710 $D=4
M629 255 63 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=51830 $Y=-10960 $D=4
M630 VDD 79 249 VDD PM L=1.8e-07 W=8.8e-07 $X=52130 $Y=-39660 $D=4
M631 VDD 80 250 VDD PM L=1.8e-07 W=8.8e-07 $X=52130 $Y=1990 $D=4
M632 263 93 68 VDD PM L=1.8e-07 W=4.4e-07 $X=52730 $Y=-13320 $D=4
M633 262 90 68 VDD PM L=1.8e-07 W=4.4e-07 $X=52780 $Y=-23910 $D=4
M634 538 79 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=52850 $Y=-39660 $D=4
M635 539 80 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=52850 $Y=1990 $D=4
M636 540 75 538 VDD PM L=1.8e-07 W=8.8e-07 $X=53280 $Y=-39660 $D=4
M637 541 76 539 VDD PM L=1.8e-07 W=8.8e-07 $X=53280 $Y=1990 $D=4
M638 280 72 540 VDD PM L=1.8e-07 W=8.8e-07 $X=53710 $Y=-39660 $D=4
M639 281 73 541 VDD PM L=1.8e-07 W=8.8e-07 $X=53710 $Y=1990 $D=4
M640 266 256 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=54140 $Y=-49810 $D=4
M641 267 257 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=54140 $Y=12580 $D=4
M642 277 264 280 VDD PM L=1.8e-07 W=8.8e-07 $X=54430 $Y=-39660 $D=4
M643 278 265 281 VDD PM L=1.8e-07 W=8.8e-07 $X=54430 $Y=1990 $D=4
M644 268 260 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54490 $Y=-26710 $D=4
M645 269 261 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54490 $Y=-10960 $D=4
M646 270 252 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54530 $Y=-36860 $D=4
M647 271 253 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=54530 $Y=-810 $D=4
M648 272 93 71 VDD PM L=1.8e-07 W=4.4e-07 $X=54680 $Y=-13320 $D=4
M649 VDD 72 277 VDD PM L=1.8e-07 W=8.8e-07 $X=55150 $Y=-39660 $D=4
M650 VDD 73 278 VDD PM L=1.8e-07 W=8.8e-07 $X=55150 $Y=1990 $D=4
M651 84 77 268 VDD PM L=1.8e-07 W=4.4e-07 $X=55250 $Y=-26270 $D=4
M652 74 78 269 VDD PM L=1.8e-07 W=4.4e-07 $X=55250 $Y=-10960 $D=4
M653 84 81 270 VDD PM L=1.8e-07 W=4.4e-07 $X=55290 $Y=-36860 $D=4
M654 74 82 271 VDD PM L=1.8e-07 W=4.4e-07 $X=55290 $Y=-370 $D=4
M655 VDD 262 273 VDD PM L=1.8e-07 W=8.8e-07 $X=55480 $Y=-23910 $D=4
M656 277 75 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=55870 $Y=-39660 $D=4
M657 278 76 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=55870 $Y=1990 $D=4
M658 263 74 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=56200 $Y=-13320 $D=4
M659 VDD 79 277 VDD PM L=1.8e-07 W=8.8e-07 $X=56590 $Y=-39660 $D=4
M660 VDD 80 278 VDD PM L=1.8e-07 W=8.8e-07 $X=56590 $Y=1990 $D=4
M661 VDD 84 263 VDD PM L=1.8e-07 W=4.4e-07 $X=56920 $Y=-13320 $D=4
M662 86 280 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=57310 $Y=-39660 $D=4
M663 87 281 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=57310 $Y=1990 $D=4
M664 282 286 77 VDD PM L=1.8e-07 W=4.4e-07 $X=57390 $Y=-26270 $D=4
M665 VDD 84 292 VDD PM L=1.8e-07 W=8.8e-07 $X=58570 $Y=-23910 $D=4
M666 290 263 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=58860 $Y=-13320 $D=4
M667 VDD 320 88 VDD PM L=1.8e-07 W=8.8e-07 $X=59250 $Y=-39660 $D=4
M668 VDD 321 89 VDD PM L=1.8e-07 W=8.8e-07 $X=59250 $Y=1990 $D=4
M669 291 288 81 VDD PM L=1.8e-07 W=4.4e-07 $X=59290 $Y=-36860 $D=4
M670 292 74 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=59290 $Y=-23910 $D=4
M671 293 289 82 VDD PM L=1.8e-07 W=4.4e-07 $X=59290 $Y=-370 $D=4
M672 294 286 81 VDD PM L=1.8e-07 W=4.4e-07 $X=59330 $Y=-26270 $D=4
M673 295 287 82 VDD PM L=1.8e-07 W=4.4e-07 $X=59330 $Y=-10960 $D=4
M674 297 262 292 VDD PM L=1.8e-07 W=8.8e-07 $X=60010 $Y=-23910 $D=4
M675 298 83 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=60050 $Y=-49810 $D=4
M676 299 85 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=60050 $Y=12580 $D=4
M677 VDD 282 294 VDD PM L=1.8e-07 W=8.8e-07 $X=60090 $Y=-26710 $D=4
M678 VDD 283 295 VDD PM L=1.8e-07 W=8.8e-07 $X=60090 $Y=-10960 $D=4
M679 284 86 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=60810 $Y=-36860 $D=4
M680 542 89 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=60810 $Y=-10960 $D=4
M681 285 87 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=60810 $Y=-370 $D=4
M682 VDD 96 305 VDD PM L=1.8e-07 W=8.8e-07 $X=61190 $Y=-39660 $D=4
M683 VDD 97 306 VDD PM L=1.8e-07 W=8.8e-07 $X=61190 $Y=1990 $D=4
M684 543 96 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61910 $Y=-39660 $D=4
M685 544 97 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61910 $Y=1990 $D=4
M686 300 297 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61950 $Y=-23910 $D=4
M687 301 290 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=61990 $Y=-13760 $D=4
M688 320 98 543 VDD PM L=1.8e-07 W=8.8e-07 $X=62340 $Y=-39660 $D=4
M689 321 99 544 VDD PM L=1.8e-07 W=8.8e-07 $X=62340 $Y=1990 $D=4
M690 302 298 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=62710 $Y=-49810 $D=4
M691 Q5I 90 300 VDD PM L=1.8e-07 W=4.4e-07 $X=62710 $Y=-23910 $D=4
M692 303 299 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=62710 $Y=12580 $D=4
M693 Q5I 93 301 VDD PM L=1.8e-07 W=4.4e-07 $X=62750 $Y=-13320 $D=4
M694 305 94 320 VDD PM L=1.8e-07 W=8.8e-07 $X=63060 $Y=-39660 $D=4
M695 306 95 321 VDD PM L=1.8e-07 W=8.8e-07 $X=63060 $Y=1990 $D=4
M696 308 284 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=63470 $Y=-36860 $D=4
M697 309 285 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=63470 $Y=-370 $D=4
M698 VDD 98 305 VDD PM L=1.8e-07 W=8.8e-07 $X=63780 $Y=-39660 $D=4
M699 VDD 99 306 VDD PM L=1.8e-07 W=8.8e-07 $X=63780 $Y=1990 $D=4
M700 312 86 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=63900 $Y=-26710 $D=4
M701 313 87 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=63900 $Y=-10960 $D=4
M702 545 98 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=64500 $Y=-39660 $D=4
M703 546 99 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=64500 $Y=1990 $D=4
M704 316 282 312 VDD PM L=1.8e-07 W=8.8e-07 $X=64620 $Y=-26710 $D=4
M705 319 113 90 VDD PM L=1.8e-07 W=4.4e-07 $X=64800 $Y=-13320 $D=4
M706 547 96 545 VDD PM L=1.8e-07 W=8.8e-07 $X=64930 $Y=-39660 $D=4
M707 548 97 546 VDD PM L=1.8e-07 W=8.8e-07 $X=64930 $Y=1990 $D=4
M708 332 94 547 VDD PM L=1.8e-07 W=8.8e-07 $X=65360 $Y=-39660 $D=4
M709 333 95 548 VDD PM L=1.8e-07 W=8.8e-07 $X=65360 $Y=1990 $D=4
M710 329 320 332 VDD PM L=1.8e-07 W=8.8e-07 $X=66080 $Y=-39660 $D=4
M711 330 321 333 VDD PM L=1.8e-07 W=8.8e-07 $X=66080 $Y=1990 $D=4
M712 323 317 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=66560 $Y=-10960 $D=4
M713 326 113 93 VDD PM L=1.8e-07 W=4.4e-07 $X=66750 $Y=-13320 $D=4
M714 327 110 93 VDD PM L=1.8e-07 W=4.4e-07 $X=66790 $Y=-23910 $D=4
M715 VDD 94 329 VDD PM L=1.8e-07 W=8.8e-07 $X=66800 $Y=-39660 $D=4
M716 VDD 95 330 VDD PM L=1.8e-07 W=8.8e-07 $X=66800 $Y=1990 $D=4
M717 103 286 322 VDD PM L=1.8e-07 W=4.4e-07 $X=67320 $Y=-26270 $D=4
M718 100 287 323 VDD PM L=1.8e-07 W=4.4e-07 $X=67320 $Y=-10960 $D=4
M719 103 288 324 VDD PM L=1.8e-07 W=4.4e-07 $X=67360 $Y=-36860 $D=4
M720 100 289 325 VDD PM L=1.8e-07 W=4.4e-07 $X=67360 $Y=-370 $D=4
M721 329 96 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=67520 $Y=-39660 $D=4
M722 330 97 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=67520 $Y=1990 $D=4
M723 VDD 318 327 VDD PM L=1.8e-07 W=8.8e-07 $X=67550 $Y=-23910 $D=4
M724 VDD 356 94 VDD PM L=1.8e-07 W=8.8e-07 $X=67820 $Y=-49810 $D=4
M725 VDD 357 95 VDD PM L=1.8e-07 W=8.8e-07 $X=67820 $Y=12140 $D=4
M726 VDD 98 329 VDD PM L=1.8e-07 W=8.8e-07 $X=68240 $Y=-39660 $D=4
M727 VDD 99 330 VDD PM L=1.8e-07 W=8.8e-07 $X=68240 $Y=1990 $D=4
M728 319 100 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=68270 $Y=-13320 $D=4
M729 104 332 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=68960 $Y=-39660 $D=4
M730 105 333 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=68960 $Y=1990 $D=4
M731 342 Q3I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=69340 $Y=-26270 $D=4
M732 343 Q8I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=69340 $Y=-10960 $D=4
M733 VDD 108 338 VDD PM L=1.8e-07 W=8.8e-07 $X=69760 $Y=-49810 $D=4
M734 VDD 109 341 VDD PM L=1.8e-07 W=8.8e-07 $X=69760 $Y=12140 $D=4
M735 286 101 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=70100 $Y=-36860 $D=4
M736 287 102 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=70100 $Y=-370 $D=4
M737 549 108 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=70480 $Y=-49810 $D=4
M738 550 109 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=70480 $Y=12140 $D=4
M739 VDD 104 286 VDD PM L=1.8e-07 W=4.4e-07 $X=70820 $Y=-36860 $D=4
M740 VDD 105 287 VDD PM L=1.8e-07 W=4.4e-07 $X=70820 $Y=-370 $D=4
M741 356 38 549 VDD PM L=1.8e-07 W=8.8e-07 $X=70910 $Y=-49810 $D=4
M742 357 39 550 VDD PM L=1.8e-07 W=8.8e-07 $X=70910 $Y=12140 $D=4
M743 336 319 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=70930 $Y=-13320 $D=4
M744 551 CLK 334 VDD PM L=1.8e-07 W=8.8e-07 $X=71280 $Y=-26710 $D=4
M745 552 CLK 335 VDD PM L=1.8e-07 W=8.8e-07 $X=71280 $Y=-10960 $D=4
M746 337 100 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=71360 $Y=-23910 $D=4
M747 338 106 356 VDD PM L=1.8e-07 W=8.8e-07 $X=71630 $Y=-49810 $D=4
M748 341 107 357 VDD PM L=1.8e-07 W=8.8e-07 $X=71630 $Y=12140 $D=4
M749 346 114 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=71700 $Y=-39220 $D=4
M750 347 115 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=71700 $Y=1990 $D=4
M751 553 RST 551 VDD PM L=1.8e-07 W=8.8e-07 $X=71710 $Y=-26710 $D=4
M752 554 RST 552 VDD PM L=1.8e-07 W=8.8e-07 $X=71710 $Y=-10960 $D=4
M753 VDD 342 553 VDD PM L=1.8e-07 W=8.8e-07 $X=72140 $Y=-26710 $D=4
M754 VDD 343 554 VDD PM L=1.8e-07 W=8.8e-07 $X=72140 $Y=-10960 $D=4
M755 VDD 38 338 VDD PM L=1.8e-07 W=8.8e-07 $X=72350 $Y=-49810 $D=4
M756 VDD 39 341 VDD PM L=1.8e-07 W=8.8e-07 $X=72350 $Y=12140 $D=4
M757 348 286 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=72760 $Y=-36860 $D=4
M758 349 287 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=72760 $Y=-370 $D=4
M759 350 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=72860 $Y=-26710 $D=4
M760 351 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=72860 $Y=-10960 $D=4
M761 555 38 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=73070 $Y=-49810 $D=4
M762 556 39 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=73070 $Y=12140 $D=4
M763 557 108 555 VDD PM L=1.8e-07 W=8.8e-07 $X=73500 $Y=-49810 $D=4
M764 558 109 556 VDD PM L=1.8e-07 W=8.8e-07 $X=73500 $Y=12140 $D=4
M765 370 106 557 VDD PM L=1.8e-07 W=8.8e-07 $X=73930 $Y=-49810 $D=4
M766 371 107 558 VDD PM L=1.8e-07 W=8.8e-07 $X=73930 $Y=12140 $D=4
M767 358 346 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=74360 $Y=-39220 $D=4
M768 359 347 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=74360 $Y=1990 $D=4
M769 364 356 370 VDD PM L=1.8e-07 W=8.8e-07 $X=74650 $Y=-49810 $D=4
M770 367 357 371 VDD PM L=1.8e-07 W=8.8e-07 $X=74650 $Y=12140 $D=4
M771 Q4I 110 354 VDD PM L=1.8e-07 W=4.4e-07 $X=74780 $Y=-23910 $D=4
M772 Q4I 113 355 VDD PM L=1.8e-07 W=4.4e-07 $X=74820 $Y=-13320 $D=4
M773 VDD 106 364 VDD PM L=1.8e-07 W=8.8e-07 $X=75370 $Y=-49810 $D=4
M774 VDD 107 367 VDD PM L=1.8e-07 W=8.8e-07 $X=75370 $Y=12140 $D=4
M775 VDD 350 Q3 VDD PM L=1.8e-07 W=8.8e-07 $X=75560 $Y=-26710 $D=4
M776 VDD 351 Q8 VDD PM L=1.8e-07 W=8.8e-07 $X=75560 $Y=-10960 $D=4
M777 121 348 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=75890 $Y=-36860 $D=4
M778 118 349 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=75890 $Y=-370 $D=4
M779 364 108 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=76090 $Y=-49810 $D=4
M780 367 109 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=76090 $Y=12140 $D=4
M781 INVQ3 Q3 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=76280 $Y=-26710 $D=4
M782 INVQ8 Q8 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=76280 $Y=-10960 $D=4
M783 VDD 38 364 VDD PM L=1.8e-07 W=8.8e-07 $X=76810 $Y=-49810 $D=4
M784 VDD 39 367 VDD PM L=1.8e-07 W=8.8e-07 $X=76810 $Y=12140 $D=4
M785 111 370 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=77530 $Y=-49810 $D=4
M786 112 371 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=77530 $Y=12140 $D=4
M787 378 Q2I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=78260 $Y=-26270 $D=4
M788 379 Q7I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=78260 $Y=-10960 $D=4
M789 374 123 113 VDD PM L=1.8e-07 W=4.4e-07 $X=78820 $Y=-13320 $D=4
M790 VDD 372 375 VDD PM L=1.8e-07 W=8.8e-07 $X=79620 $Y=-23910 $D=4
M791 559 CLK 376 VDD PM L=1.8e-07 W=8.8e-07 $X=80200 $Y=-26710 $D=4
M792 560 CLK 377 VDD PM L=1.8e-07 W=8.8e-07 $X=80200 $Y=-10960 $D=4
M793 380 116 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=80270 $Y=-49810 $D=4
M794 381 117 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=80270 $Y=12580 $D=4
M795 373 118 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=80340 $Y=-13320 $D=4
M796 561 RST 559 VDD PM L=1.8e-07 W=8.8e-07 $X=80630 $Y=-26710 $D=4
M797 562 RST 560 VDD PM L=1.8e-07 W=8.8e-07 $X=80630 $Y=-10960 $D=4
M798 VDD 378 561 VDD PM L=1.8e-07 W=8.8e-07 $X=81060 $Y=-26710 $D=4
M799 VDD 379 562 VDD PM L=1.8e-07 W=8.8e-07 $X=81060 $Y=-10960 $D=4
M800 382 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=81780 $Y=-26710 $D=4
M801 383 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=81780 $Y=-10960 $D=4
M802 384 380 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=82930 $Y=-49810 $D=4
M803 385 381 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=82930 $Y=12580 $D=4
M804 386 373 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=83000 $Y=-13320 $D=4
M805 387 118 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=83430 $Y=-23910 $D=4
M806 VDD 382 Q2 VDD PM L=1.8e-07 W=8.8e-07 $X=84480 $Y=-26710 $D=4
M807 VDD 383 Q7 VDD PM L=1.8e-07 W=8.8e-07 $X=84480 $Y=-10960 $D=4
M808 INVQ2 Q2 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=85200 $Y=-26710 $D=4
M809 INVQ7 Q7 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=85200 $Y=-10960 $D=4
M810 Q3I 122 396 VDD PM L=1.8e-07 W=4.4e-07 $X=86850 $Y=-23910 $D=4
M811 Q3I 123 397 VDD PM L=1.8e-07 W=4.4e-07 $X=86890 $Y=-13320 $D=4
M812 402 Q1I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=87180 $Y=-26270 $D=4
M813 403 Q6I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=87180 $Y=-10960 $D=4
M814 563 CLK 398 VDD PM L=1.8e-07 W=8.8e-07 $X=89120 $Y=-26710 $D=4
M815 564 CLK 399 VDD PM L=1.8e-07 W=8.8e-07 $X=89120 $Y=-10960 $D=4
M816 565 RST 563 VDD PM L=1.8e-07 W=8.8e-07 $X=89550 $Y=-26710 $D=4
M817 566 RST 564 VDD PM L=1.8e-07 W=8.8e-07 $X=89550 $Y=-10960 $D=4
M818 VDD 402 565 VDD PM L=1.8e-07 W=8.8e-07 $X=89980 $Y=-26710 $D=4
M819 VDD 403 566 VDD PM L=1.8e-07 W=8.8e-07 $X=89980 $Y=-10960 $D=4
M820 406 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=90700 $Y=-26710 $D=4
M821 407 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=90700 $Y=-10960 $D=4
M822 404 127 123 VDD PM L=1.8e-07 W=4.4e-07 $X=90890 $Y=-13320 $D=4
M823 VDD 400 405 VDD PM L=1.8e-07 W=8.8e-07 $X=91690 $Y=-23910 $D=4
M824 401 124 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=92410 $Y=-13320 $D=4
M825 VDD 406 Q1 VDD PM L=1.8e-07 W=8.8e-07 $X=93400 $Y=-26710 $D=4
M826 VDD 407 Q6 VDD PM L=1.8e-07 W=8.8e-07 $X=93400 $Y=-10960 $D=4
M827 INVQ1 Q1 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=94120 $Y=-26710 $D=4
M828 INVQ6 Q6 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=94120 $Y=-10960 $D=4
M829 412 401 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=95070 $Y=-13320 $D=4
M830 413 124 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=95500 $Y=-23910 $D=4
M831 420 Q0I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=96100 $Y=-26270 $D=4
M832 421 Q5I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=96100 $Y=-10960 $D=4
M833 567 CLK 416 VDD PM L=1.8e-07 W=8.8e-07 $X=98040 $Y=-26710 $D=4
M834 568 CLK 417 VDD PM L=1.8e-07 W=8.8e-07 $X=98040 $Y=-10960 $D=4
M835 569 RST 567 VDD PM L=1.8e-07 W=8.8e-07 $X=98470 $Y=-26710 $D=4
M836 570 RST 568 VDD PM L=1.8e-07 W=8.8e-07 $X=98470 $Y=-10960 $D=4
M837 VDD 420 569 VDD PM L=1.8e-07 W=8.8e-07 $X=98900 $Y=-26710 $D=4
M838 VDD 421 570 VDD PM L=1.8e-07 W=8.8e-07 $X=98900 $Y=-10960 $D=4
M839 Q2I 126 418 VDD PM L=1.8e-07 W=4.4e-07 $X=98920 $Y=-23910 $D=4
M840 Q2I 127 419 VDD PM L=1.8e-07 W=4.4e-07 $X=98960 $Y=-13320 $D=4
M841 422 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=99620 $Y=-26710 $D=4
M842 423 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=99620 $Y=-10960 $D=4
M843 VDD 422 Q0 VDD PM L=1.8e-07 W=8.8e-07 $X=102320 $Y=-26710 $D=4
M844 VDD 423 Q5 VDD PM L=1.8e-07 W=8.8e-07 $X=102320 $Y=-10960 $D=4
M845 430 429 127 VDD PM L=1.8e-07 W=4.4e-07 $X=102960 $Y=-13320 $D=4
M846 INVQ0 Q0 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=103040 $Y=-26710 $D=4
M847 INVQ5 Q5 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=103040 $Y=-10960 $D=4
M848 VDD 424 433 VDD PM L=1.8e-07 W=8.8e-07 $X=103760 $Y=-23910 $D=4
M849 425 128 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=104480 $Y=-13320 $D=4
M850 436 Q4I VDD VDD PM L=1.8e-07 W=4.4e-07 $X=105020 $Y=-10960 $D=4
M851 571 CLK 434 VDD PM L=1.8e-07 W=8.8e-07 $X=106960 $Y=-10960 $D=4
M852 435 425 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=107140 $Y=-13320 $D=4
M853 572 RST 571 VDD PM L=1.8e-07 W=8.8e-07 $X=107390 $Y=-10960 $D=4
M854 437 128 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=107570 $Y=-23910 $D=4
M855 VDD 436 572 VDD PM L=1.8e-07 W=8.8e-07 $X=107820 $Y=-10960 $D=4
M856 440 CLK VDD VDD PM L=1.8e-07 W=8.8e-07 $X=108540 $Y=-10960 $D=4
M857 Q1I 428 441 VDD PM L=1.8e-07 W=4.4e-07 $X=110990 $Y=-23910 $D=4
M858 Q1I 429 442 VDD PM L=1.8e-07 W=4.4e-07 $X=111030 $Y=-13320 $D=4
M859 VDD 440 Q4 VDD PM L=1.8e-07 W=8.8e-07 $X=111240 $Y=-10960 $D=4
M860 INVQ4 Q4 VDD VDD PM L=1.8e-07 W=8.8e-07 $X=111960 $Y=-10960 $D=4
M861 428 132 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=113770 $Y=-13320 $D=4
M862 445 428 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=116430 $Y=-13320 $D=4
X863 VDD 12 27 23 p18_CDNS_673868691721 $T=30540 -36420 1 0 $X=29630 $Y=-38210
X864 VDD 13 20 24 p18_CDNS_673868691721 $T=30540 -370 0 0 $X=29630 $Y=-800
X865 VDD 135 Q8I 36 p18_CDNS_673868691721 $T=30760 -23470 0 180 $X=29670 $Y=-25260
X866 VDD 21 150 55 p18_CDNS_673868691721 $T=33200 -36420 1 0 $X=32290 $Y=-38210
X867 VDD 22 151 56 p18_CDNS_673868691721 $T=33200 -370 0 0 $X=32290 $Y=-800
X868 VDD 148 21 43 p18_CDNS_673868691721 $T=33430 -26270 1 180 $X=32340 $Y=-26700
X869 VDD 149 22 44 p18_CDNS_673868691721 $T=33430 -10520 0 180 $X=32340 $Y=-12310
X870 VDD 167 24 44 p18_CDNS_673868691721 $T=35370 -10520 0 180 $X=34280 $Y=-12310
X871 VDD VDD 40 152 p18_CDNS_673868691721 $T=37050 -49370 1 0 $X=36140 $Y=-51160
X872 VDD VDD 28 153 p18_CDNS_673868691721 $T=37050 -39220 0 0 $X=36140 $Y=-39650
X873 VDD VDD 29 154 p18_CDNS_673868691721 $T=37050 2430 1 0 $X=36140 $Y=640
X874 VDD VDD 41 155 p18_CDNS_673868691721 $T=37050 12580 0 0 $X=36140 $Y=12150
X875 VDD 32 VDD 188 p18_CDNS_673868691721 $T=39110 -39220 0 0 $X=38200 $Y=-39650
X876 VDD 33 VDD 189 p18_CDNS_673868691721 $T=39110 2430 1 0 $X=38200 $Y=640
X877 VDD 207 37 68 p18_CDNS_673868691721 $T=42830 -23470 0 180 $X=41740 $Y=-25260
X878 VDD 201 VDD 59 p18_CDNS_673868691721 $T=44850 -13320 0 0 $X=43940 $Y=-13750
X879 VDD VDD 62 208 p18_CDNS_673868691721 $T=45620 -39220 0 0 $X=44710 $Y=-39650
X880 VDD VDD 63 209 p18_CDNS_673868691721 $T=45620 2430 1 0 $X=44710 $Y=640
X881 VDD 241 56 78 p18_CDNS_673868691721 $T=47440 -10520 0 180 $X=46350 $Y=-12310
X882 VDD 230 VDD 69 p18_CDNS_673868691721 $T=49460 -36420 1 0 $X=48550 $Y=-38210
X883 VDD 231 VDD 70 p18_CDNS_673868691721 $T=49460 -370 0 0 $X=48550 $Y=-800
X884 VDD 273 71 90 p18_CDNS_673868691721 $T=54900 -23470 0 180 $X=53810 $Y=-25260
X885 VDD VDD 98 266 p18_CDNS_673868691721 $T=57270 -49370 1 0 $X=56360 $Y=-51160
X886 VDD VDD 99 267 p18_CDNS_673868691721 $T=57270 12580 0 0 $X=56360 $Y=12150
X887 VDD 77 284 288 p18_CDNS_673868691721 $T=57340 -36420 1 0 $X=56430 $Y=-38210
X888 VDD 78 285 289 p18_CDNS_673868691721 $T=57340 -370 0 0 $X=56430 $Y=-800
X889 VDD 283 78 287 p18_CDNS_673868691721 $T=57570 -10520 0 180 $X=56480 $Y=-12310
X890 VDD 284 VDD 88 p18_CDNS_673868691721 $T=61530 -36420 1 0 $X=60620 $Y=-38210
X891 VDD 285 VDD 89 p18_CDNS_673868691721 $T=61530 -370 0 0 $X=60620 $Y=-800
X892 VDD 318 90 110 p18_CDNS_673868691721 $T=65030 -23470 0 180 $X=63940 $Y=-25260
X893 VDD VDD 96 302 p18_CDNS_673868691721 $T=65840 -49370 1 0 $X=64930 $Y=-51160
X894 VDD VDD 97 303 p18_CDNS_673868691721 $T=65840 12580 0 0 $X=64930 $Y=12150
X895 VDD 319 VDD 103 p18_CDNS_673868691721 $T=68990 -13320 0 0 $X=68080 $Y=-13750
X896 VDD 288 VDD 286 p18_CDNS_673868691721 $T=69380 -36420 1 0 $X=68470 $Y=-38210
X897 VDD 289 VDD 287 p18_CDNS_673868691721 $T=69380 -370 0 0 $X=68470 $Y=-800
X898 VDD 110 373 123 p18_CDNS_673868691721 $T=76870 -13320 0 0 $X=75960 $Y=-13750
X899 VDD 372 110 122 p18_CDNS_673868691721 $T=77100 -23470 0 180 $X=76010 $Y=-25260
X900 VDD VDD 125 358 p18_CDNS_673868691721 $T=77490 -39220 0 0 $X=76580 $Y=-39650
X901 VDD VDD 124 359 p18_CDNS_673868691721 $T=77490 2430 1 0 $X=76580 $Y=640
X902 VDD 375 113 122 p18_CDNS_673868691721 $T=79040 -23470 0 180 $X=77950 $Y=-25260
X903 VDD 373 VDD 121 p18_CDNS_673868691721 $T=81060 -13320 0 0 $X=80150 $Y=-13750
X904 VDD VDD 131 384 p18_CDNS_673868691721 $T=86060 -49370 1 0 $X=85150 $Y=-51160
X905 VDD VDD 128 385 p18_CDNS_673868691721 $T=86060 12580 0 0 $X=85150 $Y=12150
X906 VDD 122 401 127 p18_CDNS_673868691721 $T=88940 -13320 0 0 $X=88030 $Y=-13750
X907 VDD 400 122 126 p18_CDNS_673868691721 $T=89170 -23470 0 180 $X=88080 $Y=-25260
X908 VDD 405 123 126 p18_CDNS_673868691721 $T=91110 -23470 0 180 $X=90020 $Y=-25260
X909 VDD 401 VDD 125 p18_CDNS_673868691721 $T=93130 -13320 0 0 $X=92220 $Y=-13750
X910 VDD 126 425 429 p18_CDNS_673868691721 $T=101010 -13320 0 0 $X=100100 $Y=-13750
X911 VDD 424 126 428 p18_CDNS_673868691721 $T=101240 -23470 0 180 $X=100150 $Y=-25260
X912 VDD 433 127 428 p18_CDNS_673868691721 $T=103180 -23470 0 180 $X=102090 $Y=-25260
X913 VDD 425 VDD 131 p18_CDNS_673868691721 $T=105200 -13320 0 0 $X=104290 $Y=-13750
X914 VDD VDD Q0I 445 p18_CDNS_673868691721 $T=119560 -13320 0 0 $X=118650 $Y=-13750
X915 VDD VDD 27 517 p18_CDNS_673868691723 $T=32060 -23030 1 0 $X=31150 $Y=-25260
X916 VDD 153 14 518 p18_CDNS_673868691723 $T=34680 -39660 0 0 $X=33770 $Y=-40090
X917 VDD 154 15 519 p18_CDNS_673868691723 $T=34680 2870 1 0 $X=33770 $Y=640
X918 VDD VDD 32 522 p18_CDNS_673868691723 $T=36670 -26710 0 0 $X=35760 $Y=-27140
X919 VDD 182 28 523 p18_CDNS_673868691723 $T=40090 -35980 1 0 $X=39180 $Y=-38210
X920 VDD 183 29 524 p18_CDNS_673868691723 $T=40090 -810 0 0 $X=39180 $Y=-1240
X921 VDD 208 34 527 p18_CDNS_673868691723 $T=43250 -39660 0 0 $X=42340 $Y=-40090
X922 VDD 209 35 528 p18_CDNS_673868691723 $T=43250 2870 1 0 $X=42340 $Y=640
X923 VDD VDD 70 535 p18_CDNS_673868691723 $T=48740 -10080 1 0 $X=47830 $Y=-12310
X924 VDD VDD 27 520 p18_CDNS_673868691728 $T=35910 -13760 0 0 $X=35355 $Y=-14190
X925 VDD 149 29 521 p18_CDNS_673868691728 $T=37100 -10080 1 0 $X=36545 $Y=-12310
X926 VDD 228 62 534 p18_CDNS_673868691728 $T=49170 -26710 0 0 $X=48615 $Y=-27140
X927 VDD 283 87 542 p18_CDNS_673868691728 $T=61240 -10080 1 0 $X=60685 $Y=-12310
X928 VDD 152 VDD 16 30 ICV_1 $T=34680 -48930 1 0 $X=33770 $Y=-51160
X929 VDD 155 VDD 17 31 ICV_1 $T=34680 12140 0 0 $X=33770 $Y=11710
X930 VDD VDD 200 59 42 ICV_1 $T=44130 -23030 1 0 $X=43220 $Y=-25260
X931 VDD 252 VDD 62 69 ICV_1 $T=52160 -35980 1 0 $X=51250 $Y=-38210
X932 VDD 253 VDD 63 70 ICV_1 $T=52160 -810 0 0 $X=51250 $Y=-1240
X933 VDD 266 VDD 60 57 ICV_1 $T=54900 -48930 1 0 $X=53990 $Y=-51160
X934 VDD 267 VDD 61 58 ICV_1 $T=54900 12140 0 0 $X=53990 $Y=11710
X935 VDD VDD 262 84 74 ICV_1 $T=56200 -23030 1 0 $X=55290 $Y=-25260
X936 VDD 290 VDD 74 84 ICV_1 $T=59620 -13760 0 0 $X=58710 $Y=-14190
X937 VDD VDD 282 88 86 ICV_1 $T=60810 -26710 0 0 $X=59900 $Y=-27140
X938 VDD 302 VDD 83 91 ICV_1 $T=63470 -48930 1 0 $X=62560 $Y=-51160
X939 VDD 303 VDD 85 92 ICV_1 $T=63470 12140 0 0 $X=62560 $Y=11710
X940 VDD 308 VDD 86 88 ICV_1 $T=64230 -35980 1 0 $X=63320 $Y=-38210
X941 VDD 309 VDD 87 89 ICV_1 $T=64230 -810 0 0 $X=63320 $Y=-1240
X942 VDD VDD 318 103 100 ICV_1 $T=68270 -23030 1 0 $X=67360 $Y=-25260
X943 VDD 336 VDD 100 103 ICV_1 $T=71690 -13760 0 0 $X=70780 $Y=-14190
X944 VDD 348 VDD 101 104 ICV_1 $T=73520 -35980 1 0 $X=72610 $Y=-38210
X945 VDD 349 VDD 102 105 ICV_1 $T=73520 -810 0 0 $X=72610 $Y=-1240
X946 VDD 358 VDD 114 111 ICV_1 $T=75120 -39660 0 0 $X=74210 $Y=-40090
X947 VDD 359 VDD 115 112 ICV_1 $T=75120 2870 1 0 $X=74210 $Y=640
X948 VDD VDD 372 121 118 ICV_1 $T=80340 -23030 1 0 $X=79430 $Y=-25260
X949 VDD 384 VDD 116 119 ICV_1 $T=83690 -48930 1 0 $X=82780 $Y=-51160
X950 VDD 385 VDD 117 120 ICV_1 $T=83690 12140 0 0 $X=82780 $Y=11710
X951 VDD 386 VDD 118 121 ICV_1 $T=83760 -13760 0 0 $X=82850 $Y=-14190
X952 VDD VDD 400 125 124 ICV_1 $T=92410 -23030 1 0 $X=91500 $Y=-25260
X953 VDD 412 VDD 124 125 ICV_1 $T=95830 -13760 0 0 $X=94920 $Y=-14190
X954 VDD VDD 424 131 128 ICV_1 $T=104480 -23030 1 0 $X=103570 $Y=-25260
X955 VDD 435 VDD 128 131 ICV_1 $T=107900 -13760 0 0 $X=106990 $Y=-14190
X956 VDD 445 VDD 132 133 ICV_1 $T=117190 -13760 0 0 $X=116280 $Y=-14190
X957 GND 12 27 21 n18_CDNS_673868691726 $T=30540 -32975 1 0 $X=29880 $Y=-33765
X958 GND 134 Q8I 36 n18_CDNS_673868691726 $T=30720 -16765 1 180 $X=29880 $Y=-18785
X959 GND 13 20 22 n18_CDNS_673868691726 $T=30540 -3815 0 0 $X=29880 $Y=-5835
X960 GND 103 324 286 n18_CDNS_673868691726 $T=67540 -32975 0 180 $X=66700 $Y=-33765
X961 GND 100 325 287 n18_CDNS_673868691726 $T=67540 -3815 1 180 $X=66700 $Y=-5835
X962 GND Q1I 442 428 n18_CDNS_673868691726 $T=111210 -16765 1 180 $X=110370 $Y=-18785
X963 GND 144 152 159 16 30 ICV_2 $T=31260 -45925 1 0 $X=30600 $Y=-46715
X964 GND 18 153 160 14 25 ICV_2 $T=31260 -42665 0 0 $X=30600 $Y=-44685
X965 GND 19 154 161 15 26 ICV_2 $T=31260 5875 1 0 $X=30600 $Y=5085
X966 GND 145 155 162 17 31 ICV_2 $T=31260 9135 0 0 $X=30600 $Y=7115
X967 GND 188 208 214 34 40 ICV_2 $T=39830 -42665 0 0 $X=39170 $Y=-44685
X968 GND 189 209 215 35 41 ICV_2 $T=39830 5875 1 0 $X=39170 $Y=5085
X969 GND 256 266 274 60 57 ICV_2 $T=51480 -45925 1 0 $X=50820 $Y=-46715
X970 GND 257 267 275 61 58 ICV_2 $T=51480 9135 0 0 $X=50820 $Y=7115
X971 GND 298 302 310 83 91 ICV_2 $T=60050 -45925 1 0 $X=59390 $Y=-46715
X972 GND 299 303 311 85 92 ICV_2 $T=60050 9135 0 0 $X=59390 $Y=7115
X973 GND 286 348 352 101 104 ICV_2 $T=70100 -32975 1 0 $X=69440 $Y=-33765
X974 GND 287 349 353 102 105 ICV_2 $T=70100 -3815 0 0 $X=69440 $Y=-5835
X975 GND 346 358 362 114 111 ICV_2 $T=71700 -42665 0 0 $X=71040 $Y=-44685
X976 GND 347 359 363 115 112 ICV_2 $T=71700 5875 1 0 $X=71040 $Y=5085
X977 GND 380 384 390 116 119 ICV_2 $T=80270 -45925 1 0 $X=79610 $Y=-46715
X978 GND 381 385 391 117 120 ICV_2 $T=80270 9135 0 0 $X=79610 $Y=7115
X979 GND 428 445 446 132 133 ICV_2 $T=113770 -16765 0 0 $X=113110 $Y=-18785
X980 VDD 14 144 30 ICV_3 $T=30540 -49370 1 0 $X=29630 $Y=-51160
X981 VDD 12 18 25 ICV_3 $T=30540 -39220 0 0 $X=29630 $Y=-39650
X982 VDD 13 19 26 ICV_3 $T=30540 2430 1 0 $X=29630 $Y=640
X983 VDD 15 145 31 ICV_3 $T=30540 12580 0 0 $X=29630 $Y=12150
X984 VDD 79 256 57 ICV_3 $T=50760 -49370 1 0 $X=49850 $Y=-51160
X985 VDD 80 257 58 ICV_3 $T=50760 12580 0 0 $X=49850 $Y=12150
X986 VDD 75 298 91 ICV_3 $T=59330 -49370 1 0 $X=58420 $Y=-51160
X987 VDD 76 299 92 ICV_3 $T=59330 12580 0 0 $X=58420 $Y=12150
X988 VDD 101 346 111 ICV_3 $T=70980 -39220 0 0 $X=70070 $Y=-39650
X989 VDD 102 347 112 ICV_3 $T=70980 2430 1 0 $X=70070 $Y=640
X990 VDD 114 380 119 ICV_3 $T=79550 -49370 1 0 $X=78640 $Y=-51160
X991 VDD 115 381 120 ICV_3 $T=79550 12580 0 0 $X=78640 $Y=12150
X992 VDD 429 428 133 ICV_3 $T=113050 -13320 0 0 $X=112140 $Y=-13750
X993 VDD 134 VDD 147 p18_CDNS_6738686917210 $T=31300 -13760 0 0 $X=30390 $Y=-14190
X994 VDD 164 VDD 27 p18_CDNS_6738686917210 $T=34430 -23030 1 0 $X=33520 $Y=-25260
X995 VDD 163 VDD 150 p18_CDNS_6738686917210 $T=35910 -35980 1 0 $X=35000 $Y=-38210
X996 VDD 165 VDD 151 p18_CDNS_6738686917210 $T=35910 -810 0 0 $X=35000 $Y=-1240
X997 VDD VDD 178 177 p18_CDNS_6738686917210 $T=37810 -23030 1 0 $X=36900 $Y=-25260
X998 VDD 184 198 148 p18_CDNS_6738686917210 $T=40480 -26710 0 0 $X=39570 $Y=-27140
X999 VDD 206 VDD 201 p18_CDNS_6738686917210 $T=43370 -13760 0 0 $X=42460 $Y=-14190
X1000 VDD 233 VDD 230 p18_CDNS_6738686917210 $T=47980 -35980 1 0 $X=47070 $Y=-38210
X1001 VDD 235 VDD 231 p18_CDNS_6738686917210 $T=47980 -810 0 0 $X=47070 $Y=-1240
X1002 VDD VDD 247 232 p18_CDNS_6738686917210 $T=49920 -13760 0 0 $X=49010 $Y=-14190
X1003 VDD 255 261 229 p18_CDNS_6738686917210 $T=52550 -10080 1 0 $X=51640 $Y=-12310
X1004 VDD 272 VDD 263 p18_CDNS_6738686917210 $T=55440 -13760 0 0 $X=54530 $Y=-14190
X1005 VDD 291 VDD 284 p18_CDNS_6738686917210 $T=60050 -35980 1 0 $X=59140 $Y=-38210
X1006 VDD 293 VDD 285 p18_CDNS_6738686917210 $T=60050 -810 0 0 $X=59140 $Y=-1240
X1007 VDD 312 VDD 88 p18_CDNS_6738686917210 $T=63180 -26710 0 0 $X=62270 $Y=-27140
X1008 VDD VDD 322 316 p18_CDNS_6738686917210 $T=66560 -26710 0 0 $X=65650 $Y=-27140
X1009 VDD VDD 324 308 p18_CDNS_6738686917210 $T=66600 -35980 1 0 $X=65690 $Y=-38210
X1010 VDD VDD 325 309 p18_CDNS_6738686917210 $T=66600 -810 0 0 $X=65690 $Y=-1240
X1011 VDD 326 VDD 319 p18_CDNS_6738686917210 $T=67510 -13760 0 0 $X=66600 $Y=-14190
X1012 VDD VDD 354 345 p18_CDNS_6738686917210 $T=74020 -23030 1 0 $X=73110 $Y=-25260
X1013 VDD VDD 355 336 p18_CDNS_6738686917210 $T=74060 -13760 0 0 $X=73150 $Y=-14190
X1014 VDD 374 VDD 373 p18_CDNS_6738686917210 $T=79580 -13760 0 0 $X=78670 $Y=-14190
X1015 VDD VDD 396 393 p18_CDNS_6738686917210 $T=86090 -23030 1 0 $X=85180 $Y=-25260
X1016 VDD VDD 397 386 p18_CDNS_6738686917210 $T=86130 -13760 0 0 $X=85220 $Y=-14190
X1017 VDD 404 VDD 401 p18_CDNS_6738686917210 $T=91650 -13760 0 0 $X=90740 $Y=-14190
X1018 VDD VDD 418 415 p18_CDNS_6738686917210 $T=98160 -23030 1 0 $X=97250 $Y=-25260
X1019 VDD VDD 419 412 p18_CDNS_6738686917210 $T=98200 -13760 0 0 $X=97290 $Y=-14190
X1020 VDD 430 VDD 425 p18_CDNS_6738686917210 $T=103720 -13760 0 0 $X=102810 $Y=-14190
X1021 VDD VDD 441 439 p18_CDNS_6738686917210 $T=110230 -23030 1 0 $X=109320 $Y=-25260
X1022 VDD VDD 442 435 p18_CDNS_6738686917210 $T=110270 -13760 0 0 $X=109360 $Y=-14190
X1023 VDD 185 199 33 149 ICV_4 $T=39040 -10080 1 0 $X=38130 $Y=-12310
X1024 VDD 234 245 59 200 ICV_4 $T=46500 -23030 1 0 $X=45590 $Y=-25260
X1025 VDD 254 260 69 228 ICV_4 $T=51110 -26710 0 0 $X=50200 $Y=-27140
X1026 VDD 313 317 89 283 ICV_4 $T=63180 -10080 1 0 $X=62270 $Y=-12310
X1027 VDD 337 345 103 318 ICV_4 $T=70640 -23030 1 0 $X=69730 $Y=-25260
X1028 VDD 387 393 121 372 ICV_4 $T=82710 -23030 1 0 $X=81800 $Y=-25260
X1029 VDD 413 415 125 400 ICV_4 $T=94780 -23030 1 0 $X=93870 $Y=-25260
X1030 VDD 437 439 131 424 ICV_4 $T=106850 -23030 1 0 $X=105940 $Y=-25260
X1031 GND 146 20 n18_CDNS_6738686917211 $T=32700 -20145 1 0 $X=32000 $Y=-20715
X1032 GND 148 28 n18_CDNS_6738686917211 $T=37310 -29595 0 0 $X=36610 $Y=-31735
X1033 GND 149 29 n18_CDNS_6738686917211 $T=37310 -7195 1 0 $X=36610 $Y=-7765
X1034 GND 200 42 n18_CDNS_6738686917211 $T=44770 -20145 1 0 $X=44070 $Y=-20715
X1035 GND 228 62 n18_CDNS_6738686917211 $T=49380 -29595 0 0 $X=48680 $Y=-31735
X1036 GND 229 63 n18_CDNS_6738686917211 $T=49380 -7195 1 0 $X=48680 $Y=-7765
X1037 GND 262 74 n18_CDNS_6738686917211 $T=56840 -20145 1 0 $X=56140 $Y=-20715
X1038 GND 282 86 n18_CDNS_6738686917211 $T=61450 -29595 0 0 $X=60750 $Y=-31735
X1039 GND 283 87 n18_CDNS_6738686917211 $T=61450 -7195 1 0 $X=60750 $Y=-7765
X1040 GND 318 100 n18_CDNS_6738686917211 $T=68910 -20145 1 0 $X=68210 $Y=-20715
X1041 GND 372 118 n18_CDNS_6738686917211 $T=80980 -20145 1 0 $X=80280 $Y=-20715
X1042 GND 400 124 n18_CDNS_6738686917211 $T=93050 -20145 1 0 $X=92350 $Y=-20715
X1043 GND 424 128 n18_CDNS_6738686917211 $T=105120 -20145 1 0 $X=104420 $Y=-20715
X1044 21 148 55 GND n18_CDNS_673868691729 $T=33090 -29715 0 0 $X=32430 $Y=-30065
X1045 22 149 56 GND n18_CDNS_673868691729 $T=33090 -7075 1 0 $X=32430 $Y=-7865
X1046 36 200 71 GND n18_CDNS_673868691729 $T=40550 -20025 1 0 $X=39890 $Y=-20815
X1047 43 228 81 GND n18_CDNS_673868691729 $T=45160 -29715 0 0 $X=44500 $Y=-30065
X1048 44 229 82 GND n18_CDNS_673868691729 $T=45160 -7075 1 0 $X=44500 $Y=-7865
X1049 68 262 93 GND n18_CDNS_673868691729 $T=52620 -20025 1 0 $X=51960 $Y=-20815
X1050 77 282 288 GND n18_CDNS_673868691729 $T=57230 -29715 0 0 $X=56570 $Y=-30065
X1051 78 283 289 GND n18_CDNS_673868691729 $T=57230 -7075 1 0 $X=56570 $Y=-7865
X1052 90 318 113 GND n18_CDNS_673868691729 $T=64690 -20025 1 0 $X=64030 $Y=-20815
X1053 110 372 123 GND n18_CDNS_673868691729 $T=76760 -20025 1 0 $X=76100 $Y=-20815
X1054 122 400 127 GND n18_CDNS_673868691729 $T=88830 -20025 1 0 $X=88170 $Y=-20815
X1055 126 424 429 GND n18_CDNS_673868691729 $T=100900 -20025 1 0 $X=100240 $Y=-20815
X1056 GND 163 23 150 21 43 ICV_5 $T=33380 -32975 0 180 $X=32540 $Y=-33765
X1057 GND 165 24 151 22 44 ICV_5 $T=33380 -3815 1 180 $X=32540 $Y=-5835
X1058 GND Q7I 179 206 37 201 36 68 ICV_6 $T=38790 -16765 1 180 $X=37950 $Y=-18785
X1059 GND 59 204 233 55 230 43 77 ICV_6 $T=43400 -32975 0 180 $X=42560 $Y=-33765
X1060 GND 42 205 235 56 231 44 78 ICV_6 $T=43400 -3815 1 180 $X=42560 $Y=-5835
X1061 GND Q6I 247 272 71 263 68 90 ICV_6 $T=50860 -16765 1 180 $X=50020 $Y=-18785
X1062 GND 84 270 291 81 284 77 286 ICV_6 $T=55470 -32975 0 180 $X=54630 $Y=-33765
X1063 GND 74 271 293 82 285 78 287 ICV_6 $T=55470 -3815 1 180 $X=54630 $Y=-5835
X1064 GND Q5I 301 326 93 319 90 110 ICV_6 $T=62930 -16765 1 180 $X=62090 $Y=-18785
X1065 GND Q4I 355 374 113 373 110 122 ICV_6 $T=75000 -16765 1 180 $X=74160 $Y=-18785
X1066 GND Q3I 397 404 123 401 122 126 ICV_6 $T=87070 -16765 1 180 $X=86230 $Y=-18785
X1067 GND Q2I 419 430 127 425 126 428 ICV_6 $T=99140 -16765 1 180 $X=98300 $Y=-18785
X1068 GND 137 136 A2 A3 16 25 B3 ICV_8 $T=30540 -61490 1 0 $X=29840 $Y=-62060
X1069 GND 139 138 A0 A1 83 66 B3 ICV_8 $T=30540 -54870 1 0 $X=29840 $Y=-55440
X1070 GND 141 140 Y1 Y0 67 85 X3 ICV_8 $T=30540 16500 1 0 $X=29840 $Y=15930
X1071 GND 143 142 Y3 Y2 26 17 X3 ICV_8 $T=30540 23120 1 0 $X=29840 $Y=22550
X1072 GND 169 168 A2 A3 64 30 B2 ICV_8 $T=35390 -61490 1 0 $X=34690 $Y=-62060
X1073 GND 171 170 A0 A1 108 91 B2 ICV_8 $T=35390 -54870 1 0 $X=34690 $Y=-55440
X1074 GND 173 172 Y1 Y0 92 109 X2 ICV_8 $T=35390 16500 1 0 $X=34690 $Y=15930
X1075 GND 175 174 Y3 Y2 31 65 X2 ICV_8 $T=35390 23120 1 0 $X=34690 $Y=22550
X1076 GND 191 190 A2 A3 60 53 B1 ICV_8 $T=40240 -61490 1 0 $X=39540 $Y=-62060
X1077 GND 193 192 A0 A1 116 38 B1 ICV_8 $T=40240 -54870 1 0 $X=39540 $Y=-55440
X1078 GND 195 194 Y1 Y0 39 117 X1 ICV_8 $T=40240 16500 1 0 $X=39540 $Y=15930
X1079 GND 197 196 Y3 Y2 54 61 X1 ICV_8 $T=40240 23120 1 0 $X=39540 $Y=22550
X1080 GND 221 220 A2 A3 106 57 B0 ICV_8 $T=45090 -61490 1 0 $X=44390 $Y=-62060
X1081 GND 223 222 A0 A1 132 119 B0 ICV_8 $T=45090 -54870 1 0 $X=44390 $Y=-55440
X1082 GND 225 224 Y1 Y0 120 133 X0 ICV_8 $T=45090 16500 1 0 $X=44390 $Y=15930
X1083 GND 227 226 Y3 Y2 58 107 X0 ICV_8 $T=45090 23120 1 0 $X=44390 $Y=22550
X1084 VDD 139 B3 p18_CDNS_673868691720 $T=30540 -52050 0 0 $X=29630 $Y=-52480
X1085 VDD 140 X3 p18_CDNS_673868691720 $T=30540 15260 1 0 $X=29630 $Y=13590
X1086 VDD 137 138 A2 16 A1 66 B3 ICV_9 $T=30540 -58670 0 0 $X=29630 $Y=-59100
X1087 VDD 141 142 Y1 67 Y2 17 X3 ICV_9 $T=30540 19320 0 0 $X=29630 $Y=18890
X1088 VDD 169 170 A2 64 A1 91 B2 ICV_9 $T=35390 -58670 0 0 $X=34480 $Y=-59100
X1089 VDD 173 174 Y1 92 Y2 65 X2 ICV_9 $T=35390 19320 0 0 $X=34480 $Y=18890
X1090 VDD 191 192 A2 60 A1 38 B1 ICV_9 $T=40240 -58670 0 0 $X=39330 $Y=-59100
X1091 VDD 195 196 Y1 39 Y2 61 X1 ICV_9 $T=40240 19320 0 0 $X=39330 $Y=18890
X1092 VDD 221 222 A2 106 A1 119 B0 ICV_9 $T=45090 -58670 0 0 $X=44180 $Y=-59100
X1093 VDD 225 226 Y1 120 Y2 107 X0 ICV_9 $T=45090 19320 0 0 $X=44180 $Y=18890
X1094 VDD 136 A3 25 168 30 B3 B2 ICV_11 $T=30540 -62730 1 0 $X=29630 $Y=-64400
X1095 VDD 143 Y3 26 175 31 X3 X2 ICV_11 $T=30540 25940 0 0 $X=29630 $Y=25510
X1096 VDD 190 A3 53 220 57 B1 B0 ICV_11 $T=40240 -62730 1 0 $X=39330 $Y=-64400
X1097 VDD 193 A0 116 223 132 B1 B0 ICV_11 $T=40240 -52050 0 0 $X=39330 $Y=-52480
X1098 VDD 194 Y0 117 224 133 X1 X0 ICV_11 $T=40240 15260 1 0 $X=39330 $Y=13590
X1099 VDD 197 Y3 54 227 58 X1 X0 ICV_11 $T=40240 25940 0 0 $X=39330 $Y=25510
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_673604276091 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT n18_CDNS_673604276092 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=1.76e-06 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT Wdrive GND BIT INVBIT DATA WEN VDD
** N=10 EP=6 IP=16 FDC=8
M0 GND DATA 2 GND NM L=1.8e-07 W=2.2e-07 $X=-9920 $Y=3625 $D=0
M1 5 2 GND GND NM L=1.8e-07 W=2.2e-07 $X=-9120 $Y=3625 $D=0
M2 VDD DATA 2 VDD PM L=1.8e-07 W=4.4e-07 $X=-9880 $Y=5335 $D=4
M3 5 2 VDD VDD PM L=1.8e-07 W=4.4e-07 $X=-9160 $Y=5335 $D=4
X4 GND 6 GND 2 n18_CDNS_673604276091 $T=-10530 -2525 0 0 $X=-11190 $Y=-3655
X5 GND GND 10 5 n18_CDNS_673604276091 $T=-8510 -2525 0 0 $X=-9170 $Y=-3655
X6 GND 6 BIT WEN n18_CDNS_673604276092 $T=-10530 375 0 0 $X=-11190 $Y=25
X7 GND INVBIT 10 WEN n18_CDNS_673604276092 $T=-8510 375 0 0 $X=-9170 $Y=25
.ENDS
***************************************

* SPICE NETLIST
***************************************

.SUBCKT n18_CDNS_673724517281 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 NM L=1.8e-07 W=2.2e-07 $X=0 $Y=0 $D=0
.ENDS
***************************************
.SUBCKT p18_CDNS_673724517282 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 PM L=1.8e-07 W=4.4e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673724517280 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 3 2 1 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673724517284 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 4 2 3 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT p18_CDNS_673724517283 1 2 3 4
** N=5 EP=4 IP=0 FDC=1
M0 2 3 4 1 PM L=1.8e-07 W=1.32e-06 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=8 EP=5 IP=14 FDC=3
X0 1 3 7 p18_CDNS_673724517280 $T=0 0 0 0 $X=-910 $Y=-430
X1 1 4 7 8 p18_CDNS_673724517284 $T=430 0 0 0 $X=-125 $Y=-430
X2 1 2 5 8 p18_CDNS_673724517283 $T=860 0 0 0 $X=305 $Y=-430
.ENDS
***************************************
.SUBCKT 38Decoder ADD0 ADD1 O0 ADD2 O1 O2 O3 O4 O5 O6 O7 VDD GND
** N=16 EP=13 IP=124 FDC=54
M0 O0 ADD1 GND GND NM L=1.8e-07 W=2.2e-07 $X=-2740 $Y=3040 $D=0
M1 O1 ADD1 GND GND NM L=1.8e-07 W=2.2e-07 $X=880 $Y=3040 $D=0
M2 O2 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=4500 $Y=3040 $D=0
M3 O3 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=8120 $Y=3040 $D=0
M4 O4 ADD1 GND GND NM L=1.8e-07 W=2.2e-07 $X=11740 $Y=3040 $D=0
M5 O5 ADD1 GND GND NM L=1.8e-07 W=2.2e-07 $X=15360 $Y=3040 $D=0
M6 O6 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=18980 $Y=3040 $D=0
M7 13 ADD0 GND GND NM L=1.8e-07 W=2.2e-07 $X=19360 $Y=4760 $D=0
M8 GND 10 O6 GND NM L=1.8e-07 W=2.2e-07 $X=19780 $Y=3040 $D=0
M9 GND 13 O7 GND NM L=1.8e-07 W=2.2e-07 $X=21800 $Y=3040 $D=0
M10 O7 6 GND GND NM L=1.8e-07 W=2.2e-07 $X=22600 $Y=3040 $D=0
X11 GND O0 GND ADD0 n18_CDNS_673724517281 $T=-3540 3260 1 0 $X=-4240 $Y=2690
X12 GND O0 GND ADD2 n18_CDNS_673724517281 $T=-1940 3260 1 0 $X=-2640 $Y=2690
X13 GND O1 GND 13 n18_CDNS_673724517281 $T=80 3260 1 0 $X=-620 $Y=2690
X14 GND O1 GND ADD2 n18_CDNS_673724517281 $T=1680 3260 1 0 $X=980 $Y=2690
X15 GND O2 GND ADD0 n18_CDNS_673724517281 $T=3700 3260 1 0 $X=3000 $Y=2690
X16 GND O2 GND ADD2 n18_CDNS_673724517281 $T=5300 3260 1 0 $X=4600 $Y=2690
X17 GND O3 GND 13 n18_CDNS_673724517281 $T=7320 3260 1 0 $X=6620 $Y=2690
X18 GND O3 GND ADD2 n18_CDNS_673724517281 $T=8920 3260 1 0 $X=8220 $Y=2690
X19 GND O4 GND ADD0 n18_CDNS_673724517281 $T=10940 3260 1 0 $X=10240 $Y=2690
X20 GND O4 GND 10 n18_CDNS_673724517281 $T=12540 3260 1 0 $X=11840 $Y=2690
X21 GND O5 GND 13 n18_CDNS_673724517281 $T=14560 3260 1 0 $X=13860 $Y=2690
X22 GND O5 GND 10 n18_CDNS_673724517281 $T=16160 3260 1 0 $X=15460 $Y=2690
X23 GND O6 GND ADD0 n18_CDNS_673724517281 $T=18180 3260 1 0 $X=17480 $Y=2690
X24 GND GND 6 ADD1 n18_CDNS_673724517281 $T=21380 4760 0 0 $X=20680 $Y=3620
X25 GND O7 GND 10 n18_CDNS_673724517281 $T=23400 3260 1 0 $X=22700 $Y=2690
X26 GND GND 10 ADD2 n18_CDNS_673724517281 $T=23400 4760 0 0 $X=22700 $Y=3620
X27 VDD 13 ADD0 p18_CDNS_673724517282 $T=19360 8295 0 0 $X=18450 $Y=7865
X28 VDD 6 ADD1 p18_CDNS_673724517282 $T=21380 8295 0 0 $X=20470 $Y=7865
X29 VDD 10 ADD2 p18_CDNS_673724517282 $T=23400 8295 0 0 $X=22490 $Y=7865
X30 VDD O0 ADD0 ADD1 ADD2 ICV_1 $T=-3540 1090 1 0 $X=-4450 $Y=-1360
X31 VDD O1 13 ADD1 ADD2 ICV_1 $T=80 1090 1 0 $X=-830 $Y=-1360
X32 VDD O2 ADD0 6 ADD2 ICV_1 $T=3700 1090 1 0 $X=2790 $Y=-1360
X33 VDD O3 13 6 ADD2 ICV_1 $T=7320 1090 1 0 $X=6410 $Y=-1360
X34 VDD O4 ADD0 ADD1 10 ICV_1 $T=10940 1090 1 0 $X=10030 $Y=-1360
X35 VDD O5 13 ADD1 10 ICV_1 $T=14560 1090 1 0 $X=13650 $Y=-1360
X36 VDD O6 ADD0 6 10 ICV_1 $T=18180 1090 1 0 $X=17270 $Y=-1360
X37 VDD O7 13 6 10 ICV_1 $T=21800 1090 1 0 $X=20890 $Y=-1360
.ENDS
***************************************
